magic
tech sky130B
magscale 1 2
timestamp 1662773275
<< viali >>
rect 1501 33609 1535 33643
rect 4813 33609 4847 33643
rect 9229 33609 9263 33643
rect 14381 33609 14415 33643
rect 19257 33609 19291 33643
rect 33793 33609 33827 33643
rect 38761 33609 38795 33643
rect 43269 33609 43303 33643
rect 48605 33609 48639 33643
rect 53113 33609 53147 33643
rect 27997 33541 28031 33575
rect 28549 33541 28583 33575
rect 1685 33473 1719 33507
rect 4629 33473 4663 33507
rect 9413 33473 9447 33507
rect 14565 33473 14599 33507
rect 19441 33473 19475 33507
rect 24593 33473 24627 33507
rect 25053 33473 25087 33507
rect 30021 33473 30055 33507
rect 33609 33473 33643 33507
rect 38945 33473 38979 33507
rect 43453 33473 43487 33507
rect 48421 33473 48455 33507
rect 52929 33473 52963 33507
rect 57161 33473 57195 33507
rect 57897 33473 57931 33507
rect 30205 33337 30239 33371
rect 58081 33337 58115 33371
rect 6745 33269 6779 33303
rect 7297 33269 7331 33303
rect 24409 33269 24443 33303
rect 28641 33269 28675 33303
rect 35909 33269 35943 33303
rect 37565 33269 37599 33303
rect 57345 33269 57379 33303
rect 4537 33065 4571 33099
rect 19441 33065 19475 33099
rect 32505 33065 32539 33099
rect 37933 33065 37967 33099
rect 57529 33065 57563 33099
rect 4353 32861 4387 32895
rect 5181 32861 5215 32895
rect 5457 32861 5491 32895
rect 6193 32861 6227 32895
rect 18705 32861 18739 32895
rect 19257 32861 19291 32895
rect 22937 32861 22971 32895
rect 32321 32861 32355 32895
rect 36093 32861 36127 32895
rect 36369 32861 36403 32895
rect 37013 32861 37047 32895
rect 37749 32861 37783 32895
rect 39865 32861 39899 32895
rect 6837 32793 6871 32827
rect 37289 32793 37323 32827
rect 6377 32725 6411 32759
rect 7389 32725 7423 32759
rect 22753 32725 22787 32759
rect 23489 32725 23523 32759
rect 32965 32725 32999 32759
rect 35633 32725 35667 32759
rect 40049 32725 40083 32759
rect 52745 32725 52779 32759
rect 6561 32521 6595 32555
rect 39129 32521 39163 32555
rect 3433 32453 3467 32487
rect 5733 32453 5767 32487
rect 2053 32385 2087 32419
rect 2789 32385 2823 32419
rect 6377 32385 6411 32419
rect 37289 32385 37323 32419
rect 37933 32385 37967 32419
rect 1777 32317 1811 32351
rect 7021 32317 7055 32351
rect 7297 32317 7331 32351
rect 9045 32317 9079 32351
rect 2973 32181 3007 32215
rect 4629 32181 4663 32215
rect 9597 32181 9631 32215
rect 35725 32181 35759 32215
rect 36277 32181 36311 32215
rect 37473 32181 37507 32215
rect 38117 32181 38151 32215
rect 38577 32181 38611 32215
rect 37289 31977 37323 32011
rect 37749 31977 37783 32011
rect 8033 31841 8067 31875
rect 9505 31841 9539 31875
rect 38945 31841 38979 31875
rect 3157 31773 3191 31807
rect 5181 31773 5215 31807
rect 5457 31773 5491 31807
rect 6193 31773 6227 31807
rect 7021 31773 7055 31807
rect 7757 31773 7791 31807
rect 36093 31773 36127 31807
rect 36369 31773 36403 31807
rect 37105 31773 37139 31807
rect 37933 31773 37967 31807
rect 38669 31773 38703 31807
rect 4629 31637 4663 31671
rect 6377 31637 6411 31671
rect 6837 31637 6871 31671
rect 8953 31637 8987 31671
rect 35357 31637 35391 31671
rect 36737 31433 36771 31467
rect 37289 31433 37323 31467
rect 38945 31433 38979 31467
rect 5825 31365 5859 31399
rect 6377 31365 6411 31399
rect 4905 31297 4939 31331
rect 5641 31297 5675 31331
rect 6561 31297 6595 31331
rect 7297 31297 7331 31331
rect 35081 31297 35115 31331
rect 35817 31297 35851 31331
rect 36553 31297 36587 31331
rect 37473 31297 37507 31331
rect 38209 31297 38243 31331
rect 38485 31297 38519 31331
rect 39497 31297 39531 31331
rect 45845 31297 45879 31331
rect 46489 31297 46523 31331
rect 4629 31229 4663 31263
rect 7573 31229 7607 31263
rect 8585 31229 8619 31263
rect 35541 31229 35575 31263
rect 46029 31161 46063 31195
rect 4169 31093 4203 31127
rect 8033 31093 8067 31127
rect 2237 30889 2271 30923
rect 6377 30889 6411 30923
rect 6837 30889 6871 30923
rect 37289 30889 37323 30923
rect 37749 30889 37783 30923
rect 38945 30753 38979 30787
rect 1685 30685 1719 30719
rect 2421 30685 2455 30719
rect 3065 30685 3099 30719
rect 5181 30685 5215 30719
rect 5457 30685 5491 30719
rect 6193 30685 6227 30719
rect 7021 30685 7055 30719
rect 7757 30685 7791 30719
rect 8033 30685 8067 30719
rect 36093 30685 36127 30719
rect 36369 30685 36403 30719
rect 37105 30685 37139 30719
rect 37933 30685 37967 30719
rect 38669 30685 38703 30719
rect 1501 30549 1535 30583
rect 2881 30549 2915 30583
rect 4629 30549 4663 30583
rect 8953 30549 8987 30583
rect 35081 30549 35115 30583
rect 35541 30549 35575 30583
rect 5825 30345 5859 30379
rect 6561 30345 6595 30379
rect 37473 30345 37507 30379
rect 4905 30209 4939 30243
rect 5641 30209 5675 30243
rect 6377 30209 6411 30243
rect 14933 30209 14967 30243
rect 19533 30209 19567 30243
rect 4629 30141 4663 30175
rect 14841 30141 14875 30175
rect 36001 30073 36035 30107
rect 37933 30073 37967 30107
rect 4169 30005 4203 30039
rect 7113 30005 7147 30039
rect 7665 30005 7699 30039
rect 8125 30005 8159 30039
rect 15209 30005 15243 30039
rect 19533 30005 19567 30039
rect 37289 29801 37323 29835
rect 15025 29733 15059 29767
rect 3249 29665 3283 29699
rect 3801 29665 3835 29699
rect 7021 29665 7055 29699
rect 14565 29665 14599 29699
rect 16221 29665 16255 29699
rect 17969 29665 18003 29699
rect 20729 29665 20763 29699
rect 26893 29665 26927 29699
rect 28641 29665 28675 29699
rect 6009 29597 6043 29631
rect 14657 29597 14691 29631
rect 21005 29597 21039 29631
rect 36093 29597 36127 29631
rect 36369 29597 36403 29631
rect 37105 29597 37139 29631
rect 4077 29529 4111 29563
rect 7205 29529 7239 29563
rect 16497 29529 16531 29563
rect 18613 29529 18647 29563
rect 27169 29529 27203 29563
rect 5549 29461 5583 29495
rect 6193 29461 6227 29495
rect 8309 29461 8343 29495
rect 15761 29461 15795 29495
rect 19257 29461 19291 29495
rect 26433 29461 26467 29495
rect 29653 29461 29687 29495
rect 35541 29461 35575 29495
rect 4261 29257 4295 29291
rect 17601 29257 17635 29291
rect 24133 29257 24167 29291
rect 2053 29121 2087 29155
rect 2513 29121 2547 29155
rect 8585 29121 8619 29155
rect 17693 29121 17727 29155
rect 19993 29121 20027 29155
rect 24685 29121 24719 29155
rect 27353 29121 27387 29155
rect 36277 29121 36311 29155
rect 4997 29053 5031 29087
rect 6377 29053 6411 29087
rect 8125 29053 8159 29087
rect 19901 29053 19935 29087
rect 20821 29053 20855 29087
rect 26433 29053 26467 29087
rect 27537 29053 27571 29087
rect 28181 29053 28215 29087
rect 5365 28985 5399 29019
rect 5457 28985 5491 29019
rect 8769 28985 8803 29019
rect 36093 28985 36127 29019
rect 2770 28917 2804 28951
rect 6634 28917 6668 28951
rect 18889 28917 18923 28951
rect 24948 28917 24982 28951
rect 34805 28917 34839 28951
rect 5549 28713 5583 28747
rect 8217 28713 8251 28747
rect 18613 28713 18647 28747
rect 26801 28713 26835 28747
rect 27445 28713 27479 28747
rect 36277 28713 36311 28747
rect 5365 28645 5399 28679
rect 14289 28577 14323 28611
rect 5089 28509 5123 28543
rect 6193 28509 6227 28543
rect 6377 28509 6411 28543
rect 7021 28509 7055 28543
rect 7297 28509 7331 28543
rect 7941 28509 7975 28543
rect 14381 28509 14415 28543
rect 19257 28509 19291 28543
rect 26801 28509 26835 28543
rect 27537 28509 27571 28543
rect 35081 28509 35115 28543
rect 35357 28509 35391 28543
rect 36093 28509 36127 28543
rect 4445 28441 4479 28475
rect 4537 28373 4571 28407
rect 6561 28373 6595 28407
rect 8953 28373 8987 28407
rect 9597 28373 9631 28407
rect 14749 28373 14783 28407
rect 18061 28373 18095 28407
rect 19441 28373 19475 28407
rect 34161 28373 34195 28407
rect 2329 28169 2363 28203
rect 6377 28169 6411 28203
rect 36369 28169 36403 28203
rect 3801 28101 3835 28135
rect 8217 28101 8251 28135
rect 9137 28101 9171 28135
rect 20361 28101 20395 28135
rect 4997 28033 5031 28067
rect 6745 28033 6779 28067
rect 8033 28033 8067 28067
rect 16957 28033 16991 28067
rect 17877 28033 17911 28067
rect 20637 28033 20671 28067
rect 35449 28033 35483 28067
rect 36093 28033 36127 28067
rect 58081 28033 58115 28067
rect 1869 27965 1903 27999
rect 4077 27965 4111 27999
rect 6653 27965 6687 27999
rect 9045 27965 9079 27999
rect 10057 27965 10091 27999
rect 17785 27965 17819 27999
rect 18889 27965 18923 27999
rect 35173 27965 35207 27999
rect 18245 27897 18279 27931
rect 57897 27897 57931 27931
rect 4813 27829 4847 27863
rect 16773 27829 16807 27863
rect 34713 27829 34747 27863
rect 16024 27625 16058 27659
rect 17509 27625 17543 27659
rect 58081 27625 58115 27659
rect 4261 27557 4295 27591
rect 5365 27557 5399 27591
rect 5825 27489 5859 27523
rect 9689 27489 9723 27523
rect 15761 27489 15795 27523
rect 18337 27489 18371 27523
rect 19625 27489 19659 27523
rect 3249 27421 3283 27455
rect 5181 27421 5215 27455
rect 6009 27421 6043 27455
rect 7389 27421 7423 27455
rect 7573 27421 7607 27455
rect 9781 27421 9815 27455
rect 17969 27421 18003 27455
rect 2973 27353 3007 27387
rect 8033 27353 8067 27387
rect 8217 27353 8251 27387
rect 18153 27353 18187 27387
rect 19349 27353 19383 27387
rect 19441 27353 19475 27387
rect 1501 27285 1535 27319
rect 6469 27285 6503 27319
rect 6929 27285 6963 27319
rect 8953 27285 8987 27319
rect 15209 27285 15243 27319
rect 34989 27285 35023 27319
rect 3249 27081 3283 27115
rect 5457 27081 5491 27115
rect 18061 27081 18095 27115
rect 3893 27013 3927 27047
rect 15117 27013 15151 27047
rect 16865 27013 16899 27047
rect 3985 26945 4019 26979
rect 5089 26945 5123 26979
rect 8769 26945 8803 26979
rect 14473 26945 14507 26979
rect 15301 26945 15335 26979
rect 17877 26945 17911 26979
rect 19257 26945 19291 26979
rect 23581 26945 23615 26979
rect 4997 26877 5031 26911
rect 6377 26877 6411 26911
rect 6653 26877 6687 26911
rect 8125 26877 8159 26911
rect 14565 26877 14599 26911
rect 18705 26877 18739 26911
rect 9321 26809 9355 26843
rect 11621 26809 11655 26843
rect 13645 26809 13679 26843
rect 19441 26809 19475 26843
rect 23397 26809 23431 26843
rect 2513 26741 2547 26775
rect 8585 26741 8619 26775
rect 12357 26741 12391 26775
rect 14197 26741 14231 26775
rect 17417 26741 17451 26775
rect 19993 26741 20027 26775
rect 24225 26741 24259 26775
rect 3801 26537 3835 26571
rect 10885 26537 10919 26571
rect 17509 26537 17543 26571
rect 6193 26469 6227 26503
rect 9137 26469 9171 26503
rect 12817 26469 12851 26503
rect 18153 26469 18187 26503
rect 24777 26469 24811 26503
rect 5549 26401 5583 26435
rect 6653 26401 6687 26435
rect 8125 26401 8159 26435
rect 14657 26401 14691 26435
rect 15117 26401 15151 26435
rect 19533 26401 19567 26435
rect 22109 26401 22143 26435
rect 2421 26333 2455 26367
rect 6561 26333 6595 26367
rect 8401 26333 8435 26367
rect 8953 26333 8987 26367
rect 12633 26333 12667 26367
rect 13369 26333 13403 26367
rect 14749 26333 14783 26367
rect 15761 26333 15795 26367
rect 16589 26333 16623 26367
rect 17693 26333 17727 26367
rect 19625 26333 19659 26367
rect 20453 26333 20487 26367
rect 24961 26333 24995 26367
rect 38393 26333 38427 26367
rect 5273 26265 5307 26299
rect 12173 26265 12207 26299
rect 13461 26265 13495 26299
rect 15577 26265 15611 26299
rect 22385 26265 22419 26299
rect 38209 26265 38243 26299
rect 2329 26197 2363 26231
rect 3157 26197 3191 26231
rect 16773 26197 16807 26231
rect 19993 26197 20027 26231
rect 20637 26197 20671 26231
rect 23857 26197 23891 26231
rect 5181 25993 5215 26027
rect 5733 25993 5767 26027
rect 10977 25993 11011 26027
rect 15577 25993 15611 26027
rect 19809 25993 19843 26027
rect 22385 25993 22419 26027
rect 1685 25925 1719 25959
rect 13185 25925 13219 25959
rect 14105 25925 14139 25959
rect 30297 25925 30331 25959
rect 3709 25857 3743 25891
rect 3985 25857 4019 25891
rect 7113 25857 7147 25891
rect 7941 25857 7975 25891
rect 8585 25857 8619 25891
rect 9229 25857 9263 25891
rect 11713 25857 11747 25891
rect 13829 25857 13863 25891
rect 17141 25857 17175 25891
rect 20453 25857 20487 25891
rect 22017 25857 22051 25891
rect 23857 25857 23891 25891
rect 28641 25857 28675 25891
rect 31033 25857 31067 25891
rect 1409 25789 1443 25823
rect 7205 25789 7239 25823
rect 9505 25789 9539 25823
rect 11805 25789 11839 25823
rect 17049 25789 17083 25823
rect 18061 25789 18095 25823
rect 18337 25789 18371 25823
rect 20361 25789 20395 25823
rect 21925 25789 21959 25823
rect 12633 25721 12667 25755
rect 16129 25721 16163 25755
rect 20821 25721 20855 25755
rect 23673 25721 23707 25755
rect 3157 25653 3191 25687
rect 4445 25653 4479 25687
rect 6837 25653 6871 25687
rect 8033 25653 8067 25687
rect 8677 25653 8711 25687
rect 12081 25653 12115 25687
rect 13277 25653 13311 25687
rect 17509 25653 17543 25687
rect 28089 25653 28123 25687
rect 30941 25653 30975 25687
rect 5549 25449 5583 25483
rect 9137 25449 9171 25483
rect 10885 25449 10919 25483
rect 16957 25449 16991 25483
rect 7205 25381 7239 25415
rect 10333 25381 10367 25415
rect 14381 25381 14415 25415
rect 18061 25381 18095 25415
rect 19809 25381 19843 25415
rect 6745 25313 6779 25347
rect 7941 25313 7975 25347
rect 10057 25313 10091 25347
rect 11253 25313 11287 25347
rect 12357 25313 12391 25347
rect 12633 25313 12667 25347
rect 14841 25313 14875 25347
rect 16773 25313 16807 25347
rect 26341 25313 26375 25347
rect 29837 25313 29871 25347
rect 31861 25313 31895 25347
rect 1685 25245 1719 25279
rect 2421 25245 2455 25279
rect 3801 25245 3835 25279
rect 6837 25245 6871 25279
rect 7849 25245 7883 25279
rect 8953 25245 8987 25279
rect 9965 25245 9999 25279
rect 11161 25245 11195 25279
rect 12265 25245 12299 25279
rect 13093 25245 13127 25279
rect 14749 25245 14783 25279
rect 16037 25245 16071 25279
rect 16681 25245 16715 25279
rect 17885 25245 17919 25279
rect 18705 25245 18739 25279
rect 20361 25245 20395 25279
rect 20545 25245 20579 25279
rect 21833 25245 21867 25279
rect 22017 25245 22051 25279
rect 28733 25245 28767 25279
rect 29561 25245 29595 25279
rect 31769 25245 31803 25279
rect 34989 25245 35023 25279
rect 4077 25177 4111 25211
rect 19441 25177 19475 25211
rect 19625 25177 19659 25211
rect 22201 25177 22235 25211
rect 26617 25177 26651 25211
rect 28641 25177 28675 25211
rect 34713 25177 34747 25211
rect 1501 25109 1535 25143
rect 2237 25109 2271 25143
rect 3157 25109 3191 25143
rect 6101 25109 6135 25143
rect 8217 25109 8251 25143
rect 13185 25109 13219 25143
rect 15945 25109 15979 25143
rect 18613 25109 18647 25143
rect 21373 25109 21407 25143
rect 23029 25109 23063 25143
rect 28089 25109 28123 25143
rect 31309 25109 31343 25143
rect 5273 24905 5307 24939
rect 20913 24905 20947 24939
rect 26341 24905 26375 24939
rect 12633 24837 12667 24871
rect 3709 24769 3743 24803
rect 4813 24769 4847 24803
rect 5641 24769 5675 24803
rect 6745 24769 6779 24803
rect 8953 24769 8987 24803
rect 11621 24769 11655 24803
rect 13369 24769 13403 24803
rect 14197 24769 14231 24803
rect 15025 24769 15059 24803
rect 16129 24769 16163 24803
rect 17509 24769 17543 24803
rect 18705 24769 18739 24803
rect 18889 24769 18923 24803
rect 19533 24769 19567 24803
rect 21833 24769 21867 24803
rect 22017 24769 22051 24803
rect 23765 24769 23799 24803
rect 24501 24769 24535 24803
rect 25145 24769 25179 24803
rect 26433 24769 26467 24803
rect 27445 24769 27479 24803
rect 28457 24769 28491 24803
rect 29009 24769 29043 24803
rect 30021 24769 30055 24803
rect 30941 24769 30975 24803
rect 35909 24769 35943 24803
rect 36001 24769 36035 24803
rect 3617 24701 3651 24735
rect 5733 24701 5767 24735
rect 7021 24701 7055 24735
rect 9229 24701 9263 24735
rect 13553 24701 13587 24735
rect 15117 24701 15151 24735
rect 17601 24701 17635 24735
rect 19625 24701 19659 24735
rect 21005 24701 21039 24735
rect 21097 24701 21131 24735
rect 22477 24701 22511 24735
rect 22753 24701 22787 24735
rect 25329 24701 25363 24735
rect 31033 24701 31067 24735
rect 31585 24701 31619 24735
rect 33609 24701 33643 24735
rect 33885 24701 33919 24735
rect 37381 24701 37415 24735
rect 37657 24701 37691 24735
rect 3065 24633 3099 24667
rect 4721 24633 4755 24667
rect 14657 24633 14691 24667
rect 18889 24633 18923 24667
rect 1961 24565 1995 24599
rect 2421 24565 2455 24599
rect 4077 24565 4111 24599
rect 8493 24565 8527 24599
rect 10701 24565 10735 24599
rect 14105 24565 14139 24599
rect 16037 24565 16071 24599
rect 17233 24565 17267 24599
rect 18153 24565 18187 24599
rect 19901 24565 19935 24599
rect 20545 24565 20579 24599
rect 21925 24565 21959 24599
rect 23857 24565 23891 24599
rect 27261 24565 27295 24599
rect 28365 24565 28399 24599
rect 29193 24565 29227 24599
rect 30021 24565 30055 24599
rect 35357 24565 35391 24599
rect 39129 24565 39163 24599
rect 7205 24361 7239 24395
rect 9873 24361 9907 24395
rect 10885 24361 10919 24395
rect 15485 24361 15519 24395
rect 23305 24361 23339 24395
rect 23489 24361 23523 24395
rect 25697 24361 25731 24395
rect 28273 24361 28307 24395
rect 29009 24361 29043 24395
rect 31677 24361 31711 24395
rect 34161 24361 34195 24395
rect 39037 24361 39071 24395
rect 39957 24361 39991 24395
rect 4813 24293 4847 24327
rect 7665 24293 7699 24327
rect 12633 24293 12667 24327
rect 8125 24225 8159 24259
rect 13093 24225 13127 24259
rect 14289 24225 14323 24259
rect 14749 24225 14783 24259
rect 17325 24225 17359 24259
rect 18245 24225 18279 24259
rect 18705 24225 18739 24259
rect 22661 24225 22695 24259
rect 23581 24225 23615 24259
rect 25789 24225 25823 24259
rect 29929 24225 29963 24259
rect 30205 24225 30239 24259
rect 32689 24225 32723 24259
rect 36553 24225 36587 24259
rect 3157 24157 3191 24191
rect 3801 24157 3835 24191
rect 3985 24157 4019 24191
rect 5549 24157 5583 24191
rect 6285 24157 6319 24191
rect 8033 24157 8067 24191
rect 9229 24157 9263 24191
rect 9689 24157 9723 24191
rect 13001 24157 13035 24191
rect 14657 24157 14691 24191
rect 15301 24157 15335 24191
rect 16313 24157 16347 24191
rect 18337 24157 18371 24191
rect 21373 24157 21407 24191
rect 22569 24157 22603 24191
rect 23673 24157 23707 24191
rect 25697 24157 25731 24191
rect 26525 24157 26559 24191
rect 28825 24157 28859 24191
rect 32413 24157 32447 24191
rect 35173 24157 35207 24191
rect 35633 24157 35667 24191
rect 36461 24157 36495 24191
rect 38485 24157 38519 24191
rect 38945 24157 38979 24191
rect 39865 24157 39899 24191
rect 2881 24089 2915 24123
rect 4629 24089 4663 24123
rect 12173 24089 12207 24123
rect 19625 24089 19659 24123
rect 26801 24089 26835 24123
rect 36001 24089 36035 24123
rect 1409 24021 1443 24055
rect 3801 24021 3835 24055
rect 9045 24021 9079 24055
rect 22109 24021 22143 24055
rect 22477 24021 22511 24055
rect 24501 24021 24535 24055
rect 25053 24021 25087 24055
rect 26065 24021 26099 24055
rect 38393 24021 38427 24055
rect 47593 24021 47627 24055
rect 15209 23817 15243 23851
rect 21189 23817 21223 23851
rect 24793 23817 24827 23851
rect 30389 23817 30423 23851
rect 31125 23817 31159 23851
rect 1593 23749 1627 23783
rect 5457 23749 5491 23783
rect 5673 23749 5707 23783
rect 16957 23749 16991 23783
rect 24593 23749 24627 23783
rect 28825 23749 28859 23783
rect 33977 23749 34011 23783
rect 37565 23749 37599 23783
rect 47777 23749 47811 23783
rect 2053 23681 2087 23715
rect 3065 23681 3099 23715
rect 3341 23681 3375 23715
rect 3985 23681 4019 23715
rect 4813 23681 4847 23715
rect 6561 23681 6595 23715
rect 7021 23681 7055 23715
rect 10977 23681 11011 23715
rect 13461 23681 13495 23715
rect 13921 23681 13955 23715
rect 16773 23681 16807 23715
rect 17969 23681 18003 23715
rect 19257 23681 19291 23715
rect 21097 23681 21131 23715
rect 21281 23681 21315 23715
rect 23305 23681 23339 23715
rect 25881 23681 25915 23715
rect 27077 23681 27111 23715
rect 27997 23681 28031 23715
rect 29561 23681 29595 23715
rect 30481 23681 30515 23715
rect 31217 23681 31251 23715
rect 32137 23681 32171 23715
rect 39773 23681 39807 23715
rect 57897 23681 57931 23715
rect 3893 23613 3927 23647
rect 13185 23613 13219 23647
rect 17601 23613 17635 23647
rect 18061 23613 18095 23647
rect 19717 23613 19751 23647
rect 19993 23613 20027 23647
rect 21833 23613 21867 23647
rect 22109 23613 22143 23647
rect 23581 23613 23615 23647
rect 25605 23613 25639 23647
rect 28089 23613 28123 23647
rect 29285 23613 29319 23647
rect 29469 23613 29503 23647
rect 29653 23613 29687 23647
rect 29745 23613 29779 23647
rect 33701 23613 33735 23647
rect 37289 23613 37323 23647
rect 39037 23613 39071 23647
rect 39681 23613 39715 23647
rect 40601 23613 40635 23647
rect 47593 23613 47627 23647
rect 48605 23613 48639 23647
rect 2789 23545 2823 23579
rect 4353 23545 4387 23579
rect 4905 23545 4939 23579
rect 8309 23545 8343 23579
rect 27261 23545 27295 23579
rect 2237 23477 2271 23511
rect 3157 23477 3191 23511
rect 5641 23477 5675 23511
rect 5825 23477 5859 23511
rect 6469 23477 6503 23511
rect 9689 23477 9723 23511
rect 11713 23477 11747 23511
rect 19165 23477 19199 23511
rect 24777 23477 24811 23511
rect 24961 23477 24995 23511
rect 32229 23477 32263 23511
rect 35449 23477 35483 23511
rect 58081 23477 58115 23511
rect 8309 23273 8343 23307
rect 9873 23273 9907 23307
rect 13553 23273 13587 23307
rect 18337 23273 18371 23307
rect 18705 23273 18739 23307
rect 19809 23273 19843 23307
rect 22201 23273 22235 23307
rect 27445 23273 27479 23307
rect 33977 23273 34011 23307
rect 36001 23273 36035 23307
rect 38209 23273 38243 23307
rect 2697 23205 2731 23239
rect 17233 23205 17267 23239
rect 20913 23205 20947 23239
rect 22661 23205 22695 23239
rect 24777 23205 24811 23239
rect 26525 23205 26559 23239
rect 28089 23205 28123 23239
rect 1593 23137 1627 23171
rect 3157 23137 3191 23171
rect 4169 23137 4203 23171
rect 6561 23137 6595 23171
rect 15853 23137 15887 23171
rect 18429 23137 18463 23171
rect 21005 23137 21039 23171
rect 25973 23137 26007 23171
rect 26709 23137 26743 23171
rect 28641 23137 28675 23171
rect 42533 23137 42567 23171
rect 43177 23137 43211 23171
rect 47961 23137 47995 23171
rect 48605 23137 48639 23171
rect 2053 23069 2087 23103
rect 3065 23069 3099 23103
rect 3893 23069 3927 23103
rect 9137 23069 9171 23103
rect 11345 23069 11379 23103
rect 11805 23069 11839 23103
rect 16497 23069 16531 23103
rect 17233 23069 17267 23103
rect 17417 23069 17451 23103
rect 18521 23069 18555 23103
rect 20637 23069 20671 23103
rect 20784 23069 20818 23103
rect 22017 23069 22051 23103
rect 23673 23069 23707 23103
rect 24593 23069 24627 23103
rect 24685 23069 24719 23103
rect 24869 23069 24903 23103
rect 25053 23069 25087 23103
rect 25697 23069 25731 23103
rect 25789 23069 25823 23103
rect 26065 23069 26099 23103
rect 26617 23069 26651 23103
rect 26893 23069 26927 23103
rect 26985 23069 27019 23103
rect 29561 23069 29595 23103
rect 29837 23069 29871 23103
rect 31125 23069 31159 23103
rect 34069 23069 34103 23103
rect 35449 23069 35483 23103
rect 36093 23069 36127 23103
rect 38117 23069 38151 23103
rect 43361 23069 43395 23103
rect 47777 23069 47811 23103
rect 6837 23001 6871 23035
rect 12081 23001 12115 23035
rect 15577 23001 15611 23035
rect 17601 23001 17635 23035
rect 18061 23001 18095 23035
rect 19717 23001 19751 23035
rect 21373 23001 21407 23035
rect 21833 23001 21867 23035
rect 22845 23001 22879 23035
rect 23489 23001 23523 23035
rect 23857 23001 23891 23035
rect 25513 23001 25547 23035
rect 28089 23001 28123 23035
rect 31401 23001 31435 23035
rect 2237 22933 2271 22967
rect 5641 22933 5675 22967
rect 9045 22933 9079 22967
rect 14105 22933 14139 22967
rect 16405 22933 16439 22967
rect 24409 22933 24443 22967
rect 28549 22933 28583 22967
rect 28825 22933 28859 22967
rect 32873 22933 32907 22967
rect 35357 22933 35391 22967
rect 46213 22933 46247 22967
rect 46673 22933 46707 22967
rect 47317 22933 47351 22967
rect 4537 22729 4571 22763
rect 13093 22729 13127 22763
rect 17417 22729 17451 22763
rect 20821 22729 20855 22763
rect 25329 22729 25363 22763
rect 26157 22729 26191 22763
rect 32965 22729 32999 22763
rect 25789 22661 25823 22695
rect 32229 22661 32263 22695
rect 35541 22661 35575 22695
rect 36369 22661 36403 22695
rect 40693 22661 40727 22695
rect 48329 22661 48363 22695
rect 2145 22593 2179 22627
rect 2697 22593 2731 22627
rect 4353 22593 4387 22627
rect 5181 22593 5215 22627
rect 5825 22593 5859 22627
rect 6745 22593 6779 22627
rect 9229 22593 9263 22627
rect 11529 22593 11563 22627
rect 12541 22591 12575 22625
rect 13185 22593 13219 22627
rect 13737 22593 13771 22627
rect 16129 22593 16163 22627
rect 16681 22593 16715 22627
rect 18889 22593 18923 22627
rect 19809 22593 19843 22627
rect 21189 22593 21223 22627
rect 23121 22593 23155 22627
rect 23305 22593 23339 22627
rect 23857 22593 23891 22627
rect 24133 22593 24167 22627
rect 24777 22593 24811 22627
rect 25053 22593 25087 22627
rect 25145 22593 25179 22627
rect 25973 22593 26007 22627
rect 26249 22593 26283 22627
rect 27261 22593 27295 22627
rect 27445 22593 27479 22627
rect 29837 22593 29871 22627
rect 32321 22593 32355 22627
rect 33057 22593 33091 22627
rect 36277 22593 36311 22627
rect 37749 22593 37783 22627
rect 38393 22593 38427 22627
rect 39313 22593 39347 22627
rect 40969 22593 41003 22627
rect 41613 22593 41647 22627
rect 44465 22593 44499 22627
rect 50537 22593 50571 22627
rect 51825 22593 51859 22627
rect 7021 22525 7055 22559
rect 8769 22525 8803 22559
rect 9505 22525 9539 22559
rect 10977 22525 11011 22559
rect 14013 22525 14047 22559
rect 21097 22525 21131 22559
rect 21833 22525 21867 22559
rect 22109 22525 22143 22559
rect 23949 22525 23983 22559
rect 24869 22525 24903 22559
rect 27169 22525 27203 22559
rect 28089 22525 28123 22559
rect 28365 22525 28399 22559
rect 30113 22525 30147 22559
rect 35817 22525 35851 22559
rect 41889 22525 41923 22559
rect 44557 22525 44591 22559
rect 45293 22525 45327 22559
rect 45569 22525 45603 22559
rect 48145 22525 48179 22559
rect 48605 22525 48639 22559
rect 3157 22457 3191 22491
rect 11713 22457 11747 22491
rect 15485 22457 15519 22491
rect 18429 22457 18463 22491
rect 24317 22457 24351 22491
rect 44833 22457 44867 22491
rect 47041 22457 47075 22491
rect 50721 22457 50755 22491
rect 4997 22389 5031 22423
rect 5733 22389 5767 22423
rect 12449 22389 12483 22423
rect 16037 22389 16071 22423
rect 16865 22389 16899 22423
rect 21189 22389 21223 22423
rect 23213 22389 23247 22423
rect 23857 22389 23891 22423
rect 27629 22389 27663 22423
rect 31585 22389 31619 22423
rect 34069 22389 34103 22423
rect 37841 22389 37875 22423
rect 38485 22389 38519 22423
rect 39221 22389 39255 22423
rect 42533 22389 42567 22423
rect 47593 22389 47627 22423
rect 52009 22389 52043 22423
rect 4721 22185 4755 22219
rect 13105 22185 13139 22219
rect 19349 22185 19383 22219
rect 22569 22185 22603 22219
rect 24593 22185 24627 22219
rect 28917 22185 28951 22219
rect 29929 22185 29963 22219
rect 37000 22185 37034 22219
rect 49617 22185 49651 22219
rect 51181 22185 51215 22219
rect 51990 22185 52024 22219
rect 2329 22117 2363 22151
rect 16405 22117 16439 22151
rect 17509 22117 17543 22151
rect 22937 22117 22971 22151
rect 23581 22117 23615 22151
rect 27813 22117 27847 22151
rect 27905 22117 27939 22151
rect 2053 22049 2087 22083
rect 3893 22049 3927 22083
rect 8401 22049 8435 22083
rect 9413 22049 9447 22083
rect 13369 22049 13403 22083
rect 15853 22049 15887 22083
rect 17049 22049 17083 22083
rect 18429 22049 18463 22083
rect 18613 22049 18647 22083
rect 19717 22049 19751 22083
rect 26268 22049 26302 22083
rect 31585 22049 31619 22083
rect 34069 22049 34103 22083
rect 38485 22049 38519 22083
rect 45477 22049 45511 22083
rect 48329 22049 48363 22083
rect 49525 22049 49559 22083
rect 50813 22049 50847 22083
rect 53481 22049 53515 22083
rect 1961 21981 1995 22015
rect 3249 21981 3283 22015
rect 3801 21981 3835 22015
rect 16313 21981 16347 22015
rect 17141 21981 17175 22015
rect 19625 21981 19659 22015
rect 20361 21981 20395 22015
rect 20545 21981 20579 22015
rect 21005 21981 21039 22015
rect 21189 21981 21223 22015
rect 22477 21981 22511 22015
rect 22753 21981 22787 22015
rect 23397 21981 23431 22015
rect 24501 21981 24535 22015
rect 24685 21981 24719 22015
rect 25605 21981 25639 22015
rect 26065 21981 26099 22015
rect 26893 21981 26927 22015
rect 27077 21981 27111 22015
rect 27721 21981 27755 22015
rect 27997 21981 28031 22015
rect 28181 21981 28215 22015
rect 28825 21981 28859 22015
rect 29009 21981 29043 22015
rect 30021 21981 30055 22015
rect 30481 21981 30515 22015
rect 31493 21981 31527 22015
rect 34161 21981 34195 22015
rect 35265 21981 35299 22015
rect 35633 21981 35667 22015
rect 36737 21981 36771 22015
rect 39221 21981 39255 22015
rect 40049 21981 40083 22015
rect 43637 21981 43671 22015
rect 44281 21981 44315 22015
rect 45385 21981 45419 22015
rect 47409 21981 47443 22015
rect 48237 21981 48271 22015
rect 49617 21981 49651 22015
rect 50905 21981 50939 22015
rect 51733 21981 51767 22015
rect 55413 21981 55447 22015
rect 6193 21913 6227 21947
rect 8125 21913 8159 21947
rect 9689 21913 9723 21947
rect 15577 21913 15611 21947
rect 20453 21913 20487 21947
rect 21649 21913 21683 21947
rect 21833 21913 21867 21947
rect 22017 21913 22051 21947
rect 26341 21913 26375 21947
rect 27537 21913 27571 21947
rect 3157 21845 3191 21879
rect 6653 21845 6687 21879
rect 11161 21845 11195 21879
rect 11621 21845 11655 21879
rect 14105 21845 14139 21879
rect 17969 21845 18003 21879
rect 18337 21845 18371 21879
rect 21097 21845 21131 21879
rect 24869 21845 24903 21879
rect 25513 21845 25547 21879
rect 26157 21845 26191 21879
rect 26985 21845 27019 21879
rect 30573 21845 30607 21879
rect 32321 21845 32355 21879
rect 36277 21845 36311 21879
rect 39037 21845 39071 21879
rect 39957 21845 39991 21879
rect 43821 21845 43855 21879
rect 44465 21845 44499 21879
rect 45017 21845 45051 21879
rect 46029 21845 46063 21879
rect 46581 21845 46615 21879
rect 47593 21845 47627 21879
rect 48605 21845 48639 21879
rect 49249 21845 49283 21879
rect 50169 21845 50203 21879
rect 55597 21845 55631 21879
rect 1869 21641 1903 21675
rect 4077 21641 4111 21675
rect 11805 21641 11839 21675
rect 14749 21641 14783 21675
rect 18429 21641 18463 21675
rect 28089 21641 28123 21675
rect 34253 21641 34287 21675
rect 36277 21641 36311 21675
rect 39773 21641 39807 21675
rect 46535 21641 46569 21675
rect 47777 21641 47811 21675
rect 50169 21641 50203 21675
rect 5549 21573 5583 21607
rect 8677 21573 8711 21607
rect 10977 21573 11011 21607
rect 17141 21573 17175 21607
rect 28641 21573 28675 21607
rect 30205 21573 30239 21607
rect 38301 21573 38335 21607
rect 40325 21573 40359 21607
rect 48697 21573 48731 21607
rect 5825 21505 5859 21539
rect 10425 21505 10459 21539
rect 11713 21505 11747 21539
rect 12357 21505 12391 21539
rect 14933 21505 14967 21539
rect 15761 21505 15795 21539
rect 18705 21505 18739 21539
rect 19441 21505 19475 21539
rect 22293 21505 22327 21539
rect 23305 21505 23339 21539
rect 25697 21505 25731 21539
rect 25881 21505 25915 21539
rect 26249 21505 26283 21539
rect 27169 21505 27203 21539
rect 27445 21505 27479 21539
rect 27997 21505 28031 21539
rect 28181 21505 28215 21539
rect 31217 21505 31251 21539
rect 32873 21505 32907 21539
rect 33517 21505 33551 21539
rect 34437 21505 34471 21539
rect 35449 21505 35483 21539
rect 36461 21505 36495 21539
rect 37289 21505 37323 21539
rect 38025 21505 38059 21539
rect 40417 21505 40451 21539
rect 41061 21505 41095 21539
rect 44281 21505 44315 21539
rect 45109 21505 45143 21539
rect 47593 21505 47627 21539
rect 47869 21505 47903 21539
rect 47961 21505 47995 21539
rect 48421 21505 48455 21539
rect 50629 21505 50663 21539
rect 53021 21505 53055 21539
rect 3341 21437 3375 21471
rect 3617 21437 3651 21471
rect 6377 21437 6411 21471
rect 6653 21437 6687 21471
rect 15393 21437 15427 21471
rect 15853 21437 15887 21471
rect 18429 21437 18463 21471
rect 18613 21437 18647 21471
rect 19349 21437 19383 21471
rect 19809 21437 19843 21471
rect 20269 21437 20303 21471
rect 20545 21437 20579 21471
rect 23581 21437 23615 21471
rect 25973 21437 26007 21471
rect 26065 21437 26099 21471
rect 26985 21437 27019 21471
rect 35725 21437 35759 21471
rect 40969 21437 41003 21471
rect 42625 21437 42659 21471
rect 44097 21437 44131 21471
rect 44741 21437 44775 21471
rect 50905 21437 50939 21471
rect 55413 21437 55447 21471
rect 55689 21437 55723 21471
rect 27261 21369 27295 21403
rect 27353 21369 27387 21403
rect 41429 21369 41463 21403
rect 8125 21301 8159 21335
rect 13645 21301 13679 21335
rect 17417 21301 17451 21335
rect 22385 21301 22419 21335
rect 25053 21301 25087 21335
rect 26433 21301 26467 21335
rect 31125 21301 31159 21335
rect 32689 21301 32723 21335
rect 33425 21301 33459 21335
rect 37381 21301 37415 21335
rect 47685 21301 47719 21335
rect 52837 21301 52871 21335
rect 57161 21301 57195 21335
rect 7941 21097 7975 21131
rect 16957 21097 16991 21131
rect 19441 21097 19475 21131
rect 20545 21097 20579 21131
rect 22109 21097 22143 21131
rect 23673 21097 23707 21131
rect 24409 21097 24443 21131
rect 27261 21097 27295 21131
rect 28181 21097 28215 21131
rect 31309 21097 31343 21131
rect 33517 21097 33551 21131
rect 36369 21097 36403 21131
rect 37841 21097 37875 21131
rect 47225 21097 47259 21131
rect 49341 21097 49375 21131
rect 50629 21097 50663 21131
rect 55781 21097 55815 21131
rect 21557 21029 21591 21063
rect 22753 21029 22787 21063
rect 26525 21029 26559 21063
rect 37197 21029 37231 21063
rect 48237 21029 48271 21063
rect 54217 21029 54251 21063
rect 11621 20961 11655 20995
rect 17969 20961 18003 20995
rect 21281 20961 21315 20995
rect 28365 20961 28399 20995
rect 28457 20961 28491 20995
rect 28641 20961 28675 20995
rect 29837 20961 29871 20995
rect 31769 20961 31803 20995
rect 32045 20961 32079 20995
rect 34069 20961 34103 20995
rect 40969 20961 41003 20995
rect 43361 20961 43395 20995
rect 43637 20961 43671 20995
rect 43821 20961 43855 20995
rect 46213 20961 46247 20995
rect 51733 20961 51767 20995
rect 54309 20961 54343 20995
rect 55413 20961 55447 20995
rect 1685 20893 1719 20927
rect 3801 20893 3835 20927
rect 4445 20893 4479 20927
rect 9413 20893 9447 20927
rect 13369 20893 13403 20927
rect 14105 20893 14139 20927
rect 15669 20893 15703 20927
rect 18061 20893 18095 20927
rect 19349 20893 19383 20927
rect 20361 20893 20395 20927
rect 20545 20893 20579 20927
rect 21189 20893 21223 20927
rect 22661 20893 22695 20927
rect 23857 20893 23891 20927
rect 24685 20893 24719 20927
rect 24777 20893 24811 20927
rect 24869 20893 24903 20927
rect 25053 20893 25087 20927
rect 25697 20893 25731 20927
rect 26341 20893 26375 20927
rect 27445 20893 27479 20927
rect 27721 20893 27755 20927
rect 28549 20893 28583 20927
rect 29561 20893 29595 20927
rect 34161 20893 34195 20927
rect 34805 20893 34839 20927
rect 34989 20893 35023 20927
rect 36553 20893 36587 20927
rect 37013 20893 37047 20927
rect 38025 20893 38059 20927
rect 39313 20893 39347 20927
rect 39957 20893 39991 20927
rect 40141 20893 40175 20927
rect 44281 20893 44315 20927
rect 45293 20893 45327 20927
rect 45937 20893 45971 20927
rect 47409 20893 47443 20927
rect 47501 20893 47535 20927
rect 47685 20893 47719 20927
rect 47777 20893 47811 20927
rect 48421 20893 48455 20927
rect 48605 20893 48639 20927
rect 48697 20893 48731 20927
rect 50169 20893 50203 20927
rect 50445 20893 50479 20927
rect 51089 20893 51123 20927
rect 51273 20893 51307 20927
rect 54033 20893 54067 20927
rect 54125 20893 54159 20927
rect 55505 20893 55539 20927
rect 56701 20893 56735 20927
rect 3249 20825 3283 20859
rect 6653 20825 6687 20859
rect 13093 20825 13127 20859
rect 35817 20825 35851 20859
rect 45017 20825 45051 20859
rect 49309 20825 49343 20859
rect 49525 20825 49559 20859
rect 50261 20825 50295 20859
rect 52009 20825 52043 20859
rect 56885 20825 56919 20859
rect 3893 20757 3927 20791
rect 5733 20757 5767 20791
rect 10701 20757 10735 20791
rect 14197 20757 14231 20791
rect 15209 20757 15243 20791
rect 18429 20757 18463 20791
rect 25697 20757 25731 20791
rect 27629 20757 27663 20791
rect 39129 20757 39163 20791
rect 44465 20757 44499 20791
rect 46673 20757 46707 20791
rect 49157 20757 49191 20791
rect 51181 20757 51215 20791
rect 53481 20757 53515 20791
rect 2973 20553 3007 20587
rect 3617 20553 3651 20587
rect 4537 20553 4571 20587
rect 6653 20553 6687 20587
rect 7297 20553 7331 20587
rect 9137 20553 9171 20587
rect 10977 20553 11011 20587
rect 14473 20553 14507 20587
rect 15025 20553 15059 20587
rect 23765 20553 23799 20587
rect 33885 20553 33919 20587
rect 39773 20553 39807 20587
rect 51825 20553 51859 20587
rect 52929 20553 52963 20587
rect 53297 20553 53331 20587
rect 54217 20553 54251 20587
rect 5825 20485 5859 20519
rect 7849 20485 7883 20519
rect 10241 20485 10275 20519
rect 13921 20485 13955 20519
rect 25697 20485 25731 20519
rect 32413 20485 32447 20519
rect 36461 20485 36495 20519
rect 37289 20485 37323 20519
rect 53021 20485 53055 20519
rect 53757 20485 53791 20519
rect 1961 20417 1995 20451
rect 2789 20417 2823 20451
rect 6561 20417 6595 20451
rect 7205 20417 7239 20451
rect 10057 20417 10091 20451
rect 10793 20417 10827 20451
rect 11529 20417 11563 20451
rect 14013 20417 14047 20451
rect 15945 20417 15979 20451
rect 17509 20417 17543 20451
rect 18521 20417 18555 20451
rect 19349 20417 19383 20451
rect 22201 20417 22235 20451
rect 25973 20417 26007 20451
rect 27629 20417 27663 20451
rect 28181 20417 28215 20451
rect 29377 20417 29411 20451
rect 32137 20417 32171 20451
rect 34529 20417 34563 20451
rect 37381 20417 37415 20451
rect 40325 20417 40359 20451
rect 41153 20417 41187 20451
rect 42441 20417 42475 20451
rect 43085 20417 43119 20451
rect 44005 20417 44039 20451
rect 44649 20417 44683 20451
rect 45661 20417 45695 20451
rect 46305 20417 46339 20451
rect 48053 20417 48087 20451
rect 51457 20417 51491 20451
rect 53113 20417 53147 20451
rect 2053 20349 2087 20383
rect 11805 20349 11839 20383
rect 16037 20349 16071 20383
rect 17417 20349 17451 20383
rect 18429 20349 18463 20383
rect 18889 20349 18923 20383
rect 19625 20349 19659 20383
rect 22109 20349 22143 20383
rect 29653 20349 29687 20383
rect 36737 20349 36771 20383
rect 38025 20349 38059 20383
rect 38301 20349 38335 20383
rect 43729 20349 43763 20383
rect 45385 20349 45419 20383
rect 50169 20349 50203 20383
rect 50445 20349 50479 20383
rect 51365 20349 51399 20383
rect 2329 20281 2363 20315
rect 34437 20281 34471 20315
rect 48237 20281 48271 20315
rect 52745 20281 52779 20315
rect 54033 20281 54067 20315
rect 13277 20213 13311 20247
rect 15577 20213 15611 20247
rect 16773 20213 16807 20247
rect 17785 20213 17819 20247
rect 21097 20213 21131 20247
rect 22569 20213 22603 20247
rect 24225 20213 24259 20247
rect 31125 20213 31159 20247
rect 34989 20213 35023 20247
rect 40325 20213 40359 20247
rect 41245 20213 41279 20247
rect 41797 20213 41831 20247
rect 42625 20213 42659 20247
rect 43269 20213 43303 20247
rect 44833 20213 44867 20247
rect 46489 20213 46523 20247
rect 48697 20213 48731 20247
rect 3065 20009 3099 20043
rect 10149 20009 10183 20043
rect 10793 20009 10827 20043
rect 18613 20009 18647 20043
rect 28917 20009 28951 20043
rect 32965 20009 32999 20043
rect 39865 20009 39899 20043
rect 42717 20009 42751 20043
rect 50169 20009 50203 20043
rect 50353 20009 50387 20043
rect 51089 20009 51123 20043
rect 53849 20009 53883 20043
rect 58081 20009 58115 20043
rect 2513 19941 2547 19975
rect 6469 19941 6503 19975
rect 20545 19941 20579 19975
rect 22201 19941 22235 19975
rect 29653 19941 29687 19975
rect 38669 19941 38703 19975
rect 42257 19941 42291 19975
rect 53941 19941 53975 19975
rect 2237 19873 2271 19907
rect 11253 19873 11287 19907
rect 16497 19873 16531 19907
rect 19441 19873 19475 19907
rect 21557 19873 21591 19907
rect 22661 19873 22695 19907
rect 32413 19873 32447 19907
rect 41337 19873 41371 19907
rect 41613 19873 41647 19907
rect 43269 19873 43303 19907
rect 45017 19873 45051 19907
rect 48973 19873 49007 19907
rect 52009 19873 52043 19907
rect 53021 19873 53055 19907
rect 54033 19873 54067 19907
rect 55413 19873 55447 19907
rect 56333 19873 56367 19907
rect 2145 19805 2179 19839
rect 3157 19805 3191 19839
rect 5917 19805 5951 19839
rect 8217 19805 8251 19839
rect 9505 19805 9539 19839
rect 9965 19805 9999 19839
rect 10609 19805 10643 19839
rect 14841 19805 14875 19839
rect 15577 19805 15611 19839
rect 15761 19805 15795 19839
rect 17141 19805 17175 19839
rect 17325 19805 17359 19839
rect 19533 19805 19567 19839
rect 20361 19805 20395 19839
rect 20545 19805 20579 19839
rect 21281 19805 21315 19839
rect 22569 19805 22603 19839
rect 23213 19805 23247 19839
rect 25605 19805 25639 19839
rect 25789 19805 25823 19839
rect 26341 19805 26375 19839
rect 26525 19805 26559 19839
rect 28825 19805 28859 19839
rect 29745 19805 29779 19839
rect 30665 19805 30699 19839
rect 32873 19805 32907 19839
rect 33701 19805 33735 19839
rect 35633 19805 35667 19839
rect 38025 19805 38059 19839
rect 38485 19805 38519 19839
rect 42073 19805 42107 19839
rect 43545 19805 43579 19839
rect 44189 19805 44223 19839
rect 45293 19805 45327 19839
rect 45937 19805 45971 19839
rect 49433 19805 49467 19839
rect 49617 19805 49651 19839
rect 50353 19805 50387 19839
rect 50445 19805 50479 19839
rect 51273 19805 51307 19839
rect 51917 19805 51951 19839
rect 52102 19805 52136 19839
rect 52193 19805 52227 19839
rect 52929 19805 52963 19839
rect 53757 19805 53791 19839
rect 55505 19805 55539 19839
rect 7941 19737 7975 19771
rect 11529 19737 11563 19771
rect 24869 19737 24903 19771
rect 25053 19737 25087 19771
rect 25697 19737 25731 19771
rect 27813 19737 27847 19771
rect 28181 19737 28215 19771
rect 30941 19737 30975 19771
rect 37749 19737 37783 19771
rect 39221 19737 39255 19771
rect 44465 19737 44499 19771
rect 46213 19737 46247 19771
rect 47133 19737 47167 19771
rect 48789 19737 48823 19771
rect 50629 19737 50663 19771
rect 56609 19737 56643 19771
rect 4629 19669 4663 19703
rect 9413 19669 9447 19703
rect 13001 19669 13035 19703
rect 13553 19669 13587 19703
rect 14565 19669 14599 19703
rect 18153 19669 18187 19703
rect 19901 19669 19935 19703
rect 23765 19669 23799 19703
rect 27353 19669 27387 19703
rect 33609 19669 33643 19703
rect 35541 19669 35575 19703
rect 36277 19669 36311 19703
rect 49525 19669 49559 19703
rect 51733 19669 51767 19703
rect 53297 19669 53331 19703
rect 55873 19669 55907 19703
rect 5273 19465 5307 19499
rect 7389 19465 7423 19499
rect 10241 19465 10275 19499
rect 10885 19465 10919 19499
rect 12449 19465 12483 19499
rect 14289 19465 14323 19499
rect 16773 19465 16807 19499
rect 18705 19465 18739 19499
rect 24777 19465 24811 19499
rect 26433 19465 26467 19499
rect 31033 19465 31067 19499
rect 40969 19465 41003 19499
rect 42533 19465 42567 19499
rect 43269 19465 43303 19499
rect 48605 19465 48639 19499
rect 51641 19465 51675 19499
rect 53205 19465 53239 19499
rect 56057 19465 56091 19499
rect 7849 19397 7883 19431
rect 21925 19397 21959 19431
rect 27261 19397 27295 19431
rect 28917 19397 28951 19431
rect 46581 19397 46615 19431
rect 2145 19329 2179 19363
rect 6561 19329 6595 19363
rect 6653 19329 6687 19363
rect 7205 19329 7239 19363
rect 10333 19329 10367 19363
rect 10977 19329 11011 19363
rect 11713 19329 11747 19363
rect 11805 19329 11839 19363
rect 12541 19329 12575 19363
rect 13001 19329 13035 19363
rect 17417 19329 17451 19363
rect 17877 19329 17911 19363
rect 17969 19329 18003 19363
rect 18521 19329 18555 19363
rect 19993 19329 20027 19363
rect 22017 19329 22051 19363
rect 22477 19329 22511 19363
rect 24869 19329 24903 19363
rect 25513 19329 25547 19363
rect 27077 19329 27111 19363
rect 31125 19329 31159 19363
rect 32137 19329 32171 19363
rect 34621 19329 34655 19363
rect 36185 19329 36219 19363
rect 37565 19329 37599 19363
rect 39221 19329 39255 19363
rect 41613 19329 41647 19363
rect 42625 19329 42659 19363
rect 43085 19329 43119 19363
rect 43729 19329 43763 19363
rect 44005 19329 44039 19363
rect 44649 19329 44683 19363
rect 45385 19329 45419 19363
rect 45661 19329 45695 19363
rect 46305 19329 46339 19363
rect 47961 19329 47995 19363
rect 48881 19329 48915 19363
rect 49341 19329 49375 19363
rect 51641 19329 51675 19363
rect 51825 19329 51859 19363
rect 52745 19329 52779 19363
rect 52837 19329 52871 19363
rect 53021 19329 53055 19363
rect 53665 19329 53699 19363
rect 53849 19329 53883 19363
rect 54309 19329 54343 19363
rect 2237 19261 2271 19295
rect 3525 19261 3559 19295
rect 3801 19261 3835 19295
rect 15577 19261 15611 19295
rect 16037 19261 16071 19295
rect 19901 19261 19935 19295
rect 22753 19261 22787 19295
rect 25421 19261 25455 19295
rect 29469 19261 29503 19295
rect 32413 19261 32447 19295
rect 34529 19261 34563 19295
rect 35449 19261 35483 19295
rect 35909 19261 35943 19295
rect 37657 19261 37691 19295
rect 38393 19261 38427 19295
rect 39497 19261 39531 19295
rect 41429 19261 41463 19295
rect 47593 19261 47627 19295
rect 48053 19261 48087 19295
rect 48605 19261 48639 19295
rect 48789 19261 48823 19295
rect 49525 19261 49559 19295
rect 51181 19261 51215 19295
rect 54585 19261 54619 19295
rect 2513 19193 2547 19227
rect 9137 19193 9171 19227
rect 19349 19193 19383 19227
rect 20361 19193 20395 19227
rect 3065 19125 3099 19159
rect 5825 19125 5859 19159
rect 17325 19125 17359 19159
rect 21189 19125 21223 19159
rect 24225 19125 24259 19159
rect 25789 19125 25823 19159
rect 30389 19125 30423 19159
rect 33885 19125 33919 19159
rect 44833 19125 44867 19159
rect 53849 19125 53883 19159
rect 9597 18921 9631 18955
rect 21097 18921 21131 18955
rect 22753 18921 22787 18955
rect 29009 18921 29043 18955
rect 38761 18921 38795 18955
rect 48605 18921 48639 18955
rect 50353 18921 50387 18955
rect 52193 18921 52227 18955
rect 53205 18921 53239 18955
rect 3157 18853 3191 18887
rect 20913 18853 20947 18887
rect 25053 18853 25087 18887
rect 29561 18853 29595 18887
rect 45385 18853 45419 18887
rect 49525 18853 49559 18887
rect 53113 18853 53147 18887
rect 2237 18785 2271 18819
rect 3985 18785 4019 18819
rect 10885 18785 10919 18819
rect 13001 18785 13035 18819
rect 14289 18785 14323 18819
rect 15117 18785 15151 18819
rect 16313 18785 16347 18819
rect 19717 18785 19751 18819
rect 22385 18785 22419 18819
rect 23857 18785 23891 18819
rect 27261 18785 27295 18819
rect 36737 18785 36771 18819
rect 37381 18785 37415 18819
rect 40141 18785 40175 18819
rect 43269 18785 43303 18819
rect 47501 18785 47535 18819
rect 48421 18785 48455 18819
rect 54769 18785 54803 18819
rect 2145 18717 2179 18751
rect 2973 18717 3007 18751
rect 4261 18717 4295 18751
rect 5917 18717 5951 18751
rect 6377 18717 6411 18751
rect 9689 18717 9723 18751
rect 10333 18717 10367 18751
rect 10977 18717 11011 18751
rect 13277 18717 13311 18751
rect 14381 18717 14415 18751
rect 16037 18717 16071 18751
rect 18337 18717 18371 18751
rect 18429 18717 18463 18751
rect 20361 18717 20395 18751
rect 21097 18717 21131 18751
rect 21189 18717 21223 18751
rect 22477 18717 22511 18751
rect 24869 18717 24903 18751
rect 25789 18717 25823 18751
rect 25973 18717 26007 18751
rect 30481 18717 30515 18751
rect 31401 18717 31435 18751
rect 33793 18717 33827 18751
rect 34713 18717 34747 18751
rect 37473 18717 37507 18751
rect 38761 18717 38795 18751
rect 39865 18717 39899 18751
rect 42441 18717 42475 18751
rect 43545 18717 43579 18751
rect 44189 18717 44223 18751
rect 47685 18717 47719 18751
rect 48329 18717 48363 18751
rect 49341 18717 49375 18751
rect 50169 18717 50203 18751
rect 52101 18717 52135 18751
rect 52285 18717 52319 18751
rect 54493 18717 54527 18751
rect 57805 18717 57839 18751
rect 6653 18649 6687 18683
rect 9045 18649 9079 18683
rect 20269 18649 20303 18683
rect 21373 18649 21407 18683
rect 27537 18649 27571 18683
rect 31953 18649 31987 18683
rect 33609 18649 33643 18683
rect 34989 18649 35023 18683
rect 38301 18649 38335 18683
rect 44465 18649 44499 18683
rect 45201 18649 45235 18683
rect 45845 18649 45879 18683
rect 52745 18649 52779 18683
rect 57621 18649 57655 18683
rect 2513 18581 2547 18615
rect 4905 18581 4939 18615
rect 5825 18581 5859 18615
rect 8125 18581 8159 18615
rect 10241 18581 10275 18615
rect 11529 18581 11563 18615
rect 17785 18581 17819 18615
rect 26801 18581 26835 18615
rect 41613 18581 41647 18615
rect 42533 18581 42567 18615
rect 50905 18581 50939 18615
rect 51457 18581 51491 18615
rect 4261 18377 4295 18411
rect 5089 18377 5123 18411
rect 5733 18377 5767 18411
rect 14657 18377 14691 18411
rect 15577 18377 15611 18411
rect 21189 18377 21223 18411
rect 27261 18377 27295 18411
rect 28089 18377 28123 18411
rect 29561 18377 29595 18411
rect 41061 18377 41095 18411
rect 10977 18309 11011 18343
rect 23949 18309 23983 18343
rect 30849 18309 30883 18343
rect 40325 18309 40359 18343
rect 48053 18309 48087 18343
rect 48237 18309 48271 18343
rect 2145 18241 2179 18275
rect 3893 18241 3927 18275
rect 5181 18241 5215 18275
rect 5641 18241 5675 18275
rect 6377 18241 6411 18275
rect 7010 18241 7044 18275
rect 11529 18241 11563 18275
rect 12265 18241 12299 18275
rect 13185 18241 13219 18275
rect 14749 18241 14783 18275
rect 16681 18241 16715 18275
rect 18981 18241 19015 18275
rect 22201 18241 22235 18275
rect 27169 18241 27203 18275
rect 27353 18241 27387 18275
rect 28181 18241 28215 18275
rect 29193 18241 29227 18275
rect 30941 18241 30975 18275
rect 31493 18241 31527 18275
rect 31585 18241 31619 18275
rect 32597 18241 32631 18275
rect 33241 18241 33275 18275
rect 34437 18241 34471 18275
rect 40969 18241 41003 18275
rect 41613 18241 41647 18275
rect 42441 18241 42475 18275
rect 42717 18241 42751 18275
rect 43361 18241 43395 18275
rect 44465 18241 44499 18275
rect 50813 18241 50847 18275
rect 51273 18241 51307 18275
rect 51457 18241 51491 18275
rect 52009 18241 52043 18275
rect 52193 18241 52227 18275
rect 53021 18241 53055 18275
rect 54585 18241 54619 18275
rect 56333 18241 56367 18275
rect 57897 18241 57931 18275
rect 2237 18173 2271 18207
rect 2881 18173 2915 18207
rect 3985 18173 4019 18207
rect 7297 18173 7331 18207
rect 16957 18173 16991 18207
rect 24409 18173 24443 18207
rect 24685 18173 24719 18207
rect 26157 18173 26191 18207
rect 27997 18173 28031 18207
rect 29285 18173 29319 18207
rect 32689 18173 32723 18207
rect 34621 18173 34655 18207
rect 34897 18173 34931 18207
rect 37841 18173 37875 18207
rect 38117 18173 38151 18207
rect 40049 18173 40083 18207
rect 40509 18173 40543 18207
rect 44557 18173 44591 18207
rect 45937 18173 45971 18207
rect 46857 18173 46891 18207
rect 47041 18173 47075 18207
rect 50537 18173 50571 18207
rect 52745 18173 52779 18207
rect 52929 18173 52963 18207
rect 53113 18173 53147 18207
rect 53205 18173 53239 18207
rect 54309 18173 54343 18207
rect 56241 18173 56275 18207
rect 9689 18105 9723 18139
rect 16037 18105 16071 18139
rect 18429 18105 18463 18139
rect 28549 18105 28583 18139
rect 44097 18105 44131 18139
rect 56701 18105 56735 18139
rect 6469 18037 6503 18071
rect 8769 18037 8803 18071
rect 11621 18037 11655 18071
rect 14105 18037 14139 18071
rect 20269 18037 20303 18071
rect 33241 18037 33275 18071
rect 33977 18037 34011 18071
rect 41797 18037 41831 18071
rect 43637 18037 43671 18071
rect 49065 18037 49099 18071
rect 51365 18037 51399 18071
rect 52101 18037 52135 18071
rect 53849 18037 53883 18071
rect 58081 18037 58115 18071
rect 3065 17833 3099 17867
rect 9045 17833 9079 17867
rect 11345 17833 11379 17867
rect 22845 17833 22879 17867
rect 26249 17833 26283 17867
rect 38301 17833 38335 17867
rect 41613 17833 41647 17867
rect 42395 17833 42429 17867
rect 50629 17833 50663 17867
rect 52469 17833 52503 17867
rect 53941 17833 53975 17867
rect 54125 17833 54159 17867
rect 58173 17833 58207 17867
rect 18613 17765 18647 17799
rect 19809 17765 19843 17799
rect 23489 17765 23523 17799
rect 2237 17697 2271 17731
rect 6837 17697 6871 17731
rect 14197 17697 14231 17731
rect 14841 17697 14875 17731
rect 15945 17697 15979 17731
rect 16221 17697 16255 17731
rect 17693 17697 17727 17731
rect 28917 17697 28951 17731
rect 33333 17697 33367 17731
rect 37657 17697 37691 17731
rect 40417 17697 40451 17731
rect 43821 17697 43855 17731
rect 47593 17697 47627 17731
rect 47869 17697 47903 17731
rect 48605 17697 48639 17731
rect 50445 17697 50479 17731
rect 55505 17697 55539 17731
rect 56425 17697 56459 17731
rect 56701 17697 56735 17731
rect 2145 17629 2179 17663
rect 3249 17629 3283 17663
rect 4813 17629 4847 17663
rect 5089 17629 5123 17663
rect 6561 17629 6595 17663
rect 9137 17629 9171 17663
rect 9597 17629 9631 17663
rect 14105 17629 14139 17663
rect 15301 17629 15335 17663
rect 18705 17629 18739 17663
rect 19901 17629 19935 17663
rect 20453 17629 20487 17663
rect 20821 17629 20855 17663
rect 22753 17629 22787 17663
rect 23397 17629 23431 17663
rect 27997 17629 28031 17663
rect 28181 17629 28215 17663
rect 31769 17629 31803 17663
rect 35265 17629 35299 17663
rect 35909 17629 35943 17663
rect 38117 17629 38151 17663
rect 40325 17629 40359 17663
rect 40969 17629 41003 17663
rect 41429 17629 41463 17663
rect 44189 17629 44223 17663
rect 45017 17629 45051 17663
rect 47501 17629 47535 17663
rect 48329 17629 48363 17663
rect 50353 17629 50387 17663
rect 51641 17629 51675 17663
rect 51825 17629 51859 17663
rect 52285 17629 52319 17663
rect 52469 17629 52503 17663
rect 52929 17629 52963 17663
rect 54125 17629 54159 17663
rect 54217 17629 54251 17663
rect 55597 17629 55631 17663
rect 5733 17561 5767 17595
rect 9873 17561 9907 17595
rect 11805 17561 11839 17595
rect 22293 17561 22327 17595
rect 24961 17561 24995 17595
rect 27445 17561 27479 17595
rect 31217 17561 31251 17595
rect 31953 17561 31987 17595
rect 36185 17561 36219 17595
rect 39129 17561 39163 17595
rect 39313 17561 39347 17595
rect 45201 17561 45235 17595
rect 46857 17561 46891 17595
rect 51733 17561 51767 17595
rect 53481 17561 53515 17595
rect 54401 17561 54435 17595
rect 1777 17493 1811 17527
rect 8309 17493 8343 17527
rect 13093 17493 13127 17527
rect 15485 17493 15519 17527
rect 24409 17493 24443 17527
rect 29653 17493 29687 17527
rect 34069 17493 34103 17527
rect 35357 17493 35391 17527
rect 53113 17493 53147 17527
rect 53205 17493 53239 17527
rect 53297 17493 53331 17527
rect 55965 17493 55999 17527
rect 4537 17289 4571 17323
rect 5641 17289 5675 17323
rect 9137 17289 9171 17323
rect 25053 17289 25087 17323
rect 25697 17289 25731 17323
rect 33977 17289 34011 17323
rect 35541 17289 35575 17323
rect 41889 17289 41923 17323
rect 47593 17289 47627 17323
rect 48605 17289 48639 17323
rect 55137 17289 55171 17323
rect 55505 17289 55539 17323
rect 57897 17289 57931 17323
rect 1961 17221 1995 17255
rect 11529 17221 11563 17255
rect 14381 17221 14415 17255
rect 18981 17221 19015 17255
rect 23581 17221 23615 17255
rect 26341 17221 26375 17255
rect 45385 17221 45419 17255
rect 52929 17221 52963 17255
rect 55965 17221 55999 17255
rect 4629 17153 4663 17187
rect 5273 17153 5307 17187
rect 6561 17153 6595 17187
rect 7849 17153 7883 17187
rect 10333 17153 10367 17187
rect 10793 17153 10827 17187
rect 16681 17153 16715 17187
rect 21833 17151 21867 17185
rect 22669 17151 22703 17185
rect 23305 17153 23339 17187
rect 25789 17153 25823 17187
rect 26249 17153 26283 17187
rect 28181 17153 28215 17187
rect 28365 17153 28399 17187
rect 30021 17153 30055 17187
rect 31493 17153 31527 17187
rect 34713 17153 34747 17187
rect 34989 17153 35023 17187
rect 36277 17153 36311 17187
rect 39497 17153 39531 17187
rect 41705 17153 41739 17187
rect 47777 17153 47811 17187
rect 47869 17153 47903 17187
rect 48053 17153 48087 17187
rect 48145 17153 48179 17187
rect 49433 17153 49467 17187
rect 51917 17153 51951 17187
rect 52193 17153 52227 17187
rect 52745 17153 52779 17187
rect 55045 17153 55079 17187
rect 55321 17153 55355 17187
rect 58081 17153 58115 17187
rect 1685 17085 1719 17119
rect 3709 17085 3743 17119
rect 5365 17085 5399 17119
rect 6653 17085 6687 17119
rect 13277 17085 13311 17119
rect 13553 17085 13587 17119
rect 16957 17085 16991 17119
rect 18429 17085 18463 17119
rect 20729 17085 20763 17119
rect 29193 17085 29227 17119
rect 29929 17085 29963 17119
rect 32229 17085 32263 17119
rect 32505 17085 32539 17119
rect 37289 17085 37323 17119
rect 37565 17085 37599 17119
rect 39773 17085 39807 17119
rect 42625 17085 42659 17119
rect 44097 17085 44131 17119
rect 44281 17085 44315 17119
rect 45201 17085 45235 17119
rect 45937 17085 45971 17119
rect 49709 17085 49743 17119
rect 52101 17085 52135 17119
rect 54217 17085 54251 17119
rect 6929 17017 6963 17051
rect 10241 17017 10275 17051
rect 21189 17017 21223 17051
rect 27629 17017 27663 17051
rect 29653 17017 29687 17051
rect 51181 17017 51215 17051
rect 57253 17017 57287 17051
rect 10885 16949 10919 16983
rect 15853 16949 15887 16983
rect 21925 16949 21959 16983
rect 22753 16949 22787 16983
rect 26985 16949 27019 16983
rect 30757 16949 30791 16983
rect 31309 16949 31343 16983
rect 36093 16949 36127 16983
rect 39037 16949 39071 16983
rect 41245 16949 41279 16983
rect 51733 16949 51767 16983
rect 51917 16949 51951 16983
rect 21649 16745 21683 16779
rect 27445 16745 27479 16779
rect 32781 16745 32815 16779
rect 33333 16745 33367 16779
rect 39221 16745 39255 16779
rect 39957 16745 39991 16779
rect 40693 16745 40727 16779
rect 47133 16745 47167 16779
rect 48513 16745 48547 16779
rect 50169 16745 50203 16779
rect 54309 16745 54343 16779
rect 28457 16677 28491 16711
rect 29009 16677 29043 16711
rect 49065 16677 49099 16711
rect 53297 16677 53331 16711
rect 3249 16609 3283 16643
rect 6285 16609 6319 16643
rect 6745 16609 6779 16643
rect 7849 16609 7883 16643
rect 8401 16609 8435 16643
rect 9505 16609 9539 16643
rect 12909 16609 12943 16643
rect 13185 16609 13219 16643
rect 17601 16609 17635 16643
rect 20821 16609 20855 16643
rect 21097 16609 21131 16643
rect 24409 16609 24443 16643
rect 24685 16609 24719 16643
rect 29561 16609 29595 16643
rect 30021 16609 30055 16643
rect 31309 16609 31343 16643
rect 36369 16609 36403 16643
rect 36645 16609 36679 16643
rect 42625 16609 42659 16643
rect 45661 16609 45695 16643
rect 49341 16609 49375 16643
rect 50629 16609 50663 16643
rect 51457 16609 51491 16643
rect 51733 16609 51767 16643
rect 55413 16609 55447 16643
rect 56425 16609 56459 16643
rect 56701 16609 56735 16643
rect 3893 16541 3927 16575
rect 3985 16541 4019 16575
rect 4629 16541 4663 16575
rect 5181 16541 5215 16575
rect 5273 16541 5307 16575
rect 6193 16541 6227 16575
rect 7573 16541 7607 16575
rect 9229 16541 9263 16575
rect 10885 16541 10919 16575
rect 14105 16541 14139 16575
rect 14933 16541 14967 16575
rect 15393 16541 15427 16575
rect 17877 16541 17911 16575
rect 18337 16541 18371 16575
rect 18429 16541 18463 16575
rect 22109 16541 22143 16575
rect 26617 16541 26651 16575
rect 27537 16541 27571 16575
rect 28733 16541 28767 16575
rect 29929 16541 29963 16575
rect 31033 16541 31067 16575
rect 34161 16541 34195 16575
rect 34805 16541 34839 16575
rect 34897 16541 34931 16575
rect 35449 16541 35483 16575
rect 35541 16541 35575 16575
rect 38577 16541 38611 16575
rect 40049 16541 40083 16575
rect 40785 16541 40819 16575
rect 43269 16541 43303 16575
rect 43729 16541 43763 16575
rect 45385 16541 45419 16575
rect 48053 16541 48087 16575
rect 48329 16541 48363 16575
rect 48973 16541 49007 16575
rect 50537 16541 50571 16575
rect 53849 16541 53883 16575
rect 53941 16541 53975 16575
rect 54125 16541 54159 16575
rect 55505 16541 55539 16575
rect 10793 16473 10827 16507
rect 14841 16473 14875 16507
rect 22385 16473 22419 16507
rect 26709 16473 26743 16507
rect 33425 16473 33459 16507
rect 38669 16473 38703 16507
rect 43085 16473 43119 16507
rect 4537 16405 4571 16439
rect 10057 16405 10091 16439
rect 11437 16405 11471 16439
rect 14289 16405 14323 16439
rect 15485 16405 15519 16439
rect 16129 16405 16163 16439
rect 19349 16405 19383 16439
rect 23857 16405 23891 16439
rect 26157 16405 26191 16439
rect 28641 16405 28675 16439
rect 28825 16405 28859 16439
rect 34069 16405 34103 16439
rect 38117 16405 38151 16439
rect 43913 16405 43947 16439
rect 48145 16405 48179 16439
rect 49065 16405 49099 16439
rect 49157 16405 49191 16439
rect 52745 16405 52779 16439
rect 52929 16405 52963 16439
rect 53021 16405 53055 16439
rect 53113 16405 53147 16439
rect 55873 16405 55907 16439
rect 58173 16405 58207 16439
rect 3433 16201 3467 16235
rect 31493 16201 31527 16235
rect 33885 16201 33919 16235
rect 37749 16201 37783 16235
rect 49249 16201 49283 16235
rect 50261 16201 50295 16235
rect 55137 16201 55171 16235
rect 4537 16133 4571 16167
rect 12265 16133 12299 16167
rect 19717 16133 19751 16167
rect 22201 16133 22235 16167
rect 23213 16133 23247 16167
rect 34897 16133 34931 16167
rect 39129 16133 39163 16167
rect 44741 16133 44775 16167
rect 44957 16133 44991 16167
rect 45569 16133 45603 16167
rect 48053 16133 48087 16167
rect 50905 16133 50939 16167
rect 51825 16133 51859 16167
rect 53849 16133 53883 16167
rect 55965 16133 55999 16167
rect 3985 16065 4019 16099
rect 4629 16065 4663 16099
rect 5457 16065 5491 16099
rect 6377 16065 6411 16099
rect 8769 16065 8803 16099
rect 14381 16065 14415 16099
rect 22385 16065 22419 16099
rect 22937 16065 22971 16099
rect 25421 16065 25455 16099
rect 27629 16065 27663 16099
rect 29009 16065 29043 16099
rect 29377 16065 29411 16099
rect 30757 16065 30791 16099
rect 31401 16065 31435 16099
rect 36001 16065 36035 16099
rect 37841 16065 37875 16099
rect 38393 16065 38427 16099
rect 38577 16065 38611 16099
rect 39037 16065 39071 16099
rect 39681 16065 39715 16099
rect 41061 16065 41095 16099
rect 45845 16065 45879 16099
rect 46489 16065 46523 16099
rect 47961 16065 47995 16099
rect 48237 16065 48271 16099
rect 48881 16065 48915 16099
rect 49065 16065 49099 16099
rect 50997 16065 51031 16099
rect 51917 16065 51951 16099
rect 52745 16065 52779 16099
rect 52837 16065 52871 16099
rect 53665 16065 53699 16099
rect 54677 16065 54711 16099
rect 54769 16065 54803 16099
rect 54953 16065 54987 16099
rect 55597 16065 55631 16099
rect 55781 16065 55815 16099
rect 57161 16065 57195 16099
rect 5365 15997 5399 16031
rect 10977 15997 11011 16031
rect 11989 15997 12023 16031
rect 17233 15997 17267 16031
rect 18705 15997 18739 16031
rect 18981 15997 19015 16031
rect 19441 15997 19475 16031
rect 21189 15997 21223 16031
rect 27721 15997 27755 16031
rect 28457 15997 28491 16031
rect 30021 15997 30055 16031
rect 32137 15997 32171 16031
rect 32413 15997 32447 16031
rect 35909 15997 35943 16031
rect 36369 15997 36403 16031
rect 40969 15997 41003 16031
rect 41889 15997 41923 16031
rect 42441 15997 42475 16031
rect 42717 15997 42751 16031
rect 46765 15997 46799 16031
rect 52101 15997 52135 16031
rect 53021 15997 53055 16031
rect 54033 15997 54067 16031
rect 57069 15997 57103 16031
rect 5825 15929 5859 15963
rect 6469 15929 6503 15963
rect 9229 15929 9263 15963
rect 13737 15929 13771 15963
rect 26065 15929 26099 15963
rect 39773 15929 39807 15963
rect 56793 15929 56827 15963
rect 7481 15861 7515 15895
rect 10713 15861 10747 15895
rect 15669 15861 15703 15895
rect 24685 15861 24719 15895
rect 25513 15861 25547 15895
rect 30665 15861 30699 15895
rect 34989 15861 35023 15895
rect 38577 15861 38611 15895
rect 44189 15861 44223 15895
rect 44925 15861 44959 15895
rect 45109 15861 45143 15895
rect 48421 15861 48455 15895
rect 48881 15861 48915 15895
rect 49709 15861 49743 15895
rect 51457 15861 51491 15895
rect 52929 15861 52963 15895
rect 9137 15657 9171 15691
rect 12357 15657 12391 15691
rect 14657 15657 14691 15691
rect 18613 15657 18647 15691
rect 19349 15657 19383 15691
rect 23857 15657 23891 15691
rect 24501 15657 24535 15691
rect 28273 15657 28307 15691
rect 36461 15657 36495 15691
rect 51181 15657 51215 15691
rect 53021 15657 53055 15691
rect 54125 15657 54159 15691
rect 58081 15657 58115 15691
rect 9781 15589 9815 15623
rect 15209 15589 15243 15623
rect 17969 15589 18003 15623
rect 27721 15589 27755 15623
rect 32137 15589 32171 15623
rect 44465 15589 44499 15623
rect 8309 15521 8343 15555
rect 16957 15521 16991 15555
rect 20085 15521 20119 15555
rect 21833 15521 21867 15555
rect 25421 15521 25455 15555
rect 25973 15521 26007 15555
rect 26249 15521 26283 15555
rect 28917 15521 28951 15555
rect 34713 15521 34747 15555
rect 38761 15521 38795 15555
rect 39037 15521 39071 15555
rect 39957 15521 39991 15555
rect 40417 15521 40451 15555
rect 41613 15521 41647 15555
rect 44189 15521 44223 15555
rect 45201 15521 45235 15555
rect 45937 15521 45971 15555
rect 48237 15521 48271 15555
rect 49157 15521 49191 15555
rect 54677 15521 54711 15555
rect 56333 15521 56367 15555
rect 56609 15521 56643 15555
rect 5365 15453 5399 15487
rect 5457 15453 5491 15487
rect 6561 15453 6595 15487
rect 6745 15453 6779 15487
rect 8401 15453 8435 15487
rect 9229 15453 9263 15487
rect 9689 15453 9723 15487
rect 10425 15453 10459 15487
rect 13369 15453 13403 15487
rect 14473 15453 14507 15487
rect 18061 15453 18095 15487
rect 18521 15453 18555 15487
rect 19809 15453 19843 15487
rect 22385 15453 22419 15487
rect 23029 15453 23063 15487
rect 23673 15453 23707 15487
rect 24593 15453 24627 15487
rect 25513 15453 25547 15487
rect 28181 15453 28215 15487
rect 29009 15453 29043 15487
rect 29561 15453 29595 15487
rect 33149 15453 33183 15487
rect 33333 15453 33367 15487
rect 33885 15453 33919 15487
rect 33977 15453 34011 15487
rect 37105 15453 37139 15487
rect 37657 15453 37691 15487
rect 39129 15453 39163 15487
rect 40049 15453 40083 15487
rect 40877 15453 40911 15487
rect 44097 15453 44131 15487
rect 45017 15453 45051 15487
rect 48407 15453 48441 15487
rect 50169 15453 50203 15487
rect 51089 15453 51123 15487
rect 51273 15453 51307 15487
rect 51917 15453 51951 15487
rect 52193 15453 52227 15487
rect 53941 15453 53975 15487
rect 54033 15453 54067 15487
rect 54217 15453 54251 15487
rect 11069 15385 11103 15419
rect 16681 15385 16715 15419
rect 22477 15385 22511 15419
rect 29745 15385 29779 15419
rect 31401 15385 31435 15419
rect 34989 15385 35023 15419
rect 41889 15385 41923 15419
rect 47501 15385 47535 15419
rect 49341 15385 49375 15419
rect 52101 15385 52135 15419
rect 52989 15385 53023 15419
rect 53205 15385 53239 15419
rect 6009 15317 6043 15351
rect 7573 15317 7607 15351
rect 10609 15317 10643 15351
rect 13461 15317 13495 15351
rect 23213 15317 23247 15351
rect 33241 15317 33275 15351
rect 37013 15317 37047 15351
rect 37749 15317 37783 15351
rect 40969 15317 41003 15351
rect 43361 15317 43395 15351
rect 47593 15317 47627 15351
rect 48697 15317 48731 15351
rect 50353 15317 50387 15351
rect 51733 15317 51767 15351
rect 52837 15317 52871 15351
rect 5273 15113 5307 15147
rect 15669 15113 15703 15147
rect 21281 15113 21315 15147
rect 27445 15113 27479 15147
rect 31217 15113 31251 15147
rect 32781 15113 32815 15147
rect 35357 15113 35391 15147
rect 36001 15113 36035 15147
rect 39589 15113 39623 15147
rect 40141 15113 40175 15147
rect 50721 15113 50755 15147
rect 52745 15113 52779 15147
rect 55137 15113 55171 15147
rect 8677 15045 8711 15079
rect 10701 15045 10735 15079
rect 14381 15045 14415 15079
rect 16865 15045 16899 15079
rect 21833 15045 21867 15079
rect 24685 15045 24719 15079
rect 30573 15045 30607 15079
rect 38761 15045 38795 15079
rect 42441 15045 42475 15079
rect 49249 15045 49283 15079
rect 5733 14977 5767 15011
rect 6653 14977 6687 15011
rect 7481 14977 7515 15011
rect 7941 14977 7975 15011
rect 8585 14977 8619 15011
rect 11529 14977 11563 15011
rect 16773 14977 16807 15011
rect 20637 14977 20671 15011
rect 20913 14977 20947 15011
rect 24041 14977 24075 15011
rect 27353 14977 27387 15011
rect 27997 14977 28031 15011
rect 32321 14977 32355 15011
rect 33609 14977 33643 15011
rect 36093 14977 36127 15011
rect 36737 14977 36771 15011
rect 39037 14977 39071 15011
rect 39681 14977 39715 15011
rect 40969 14977 41003 15011
rect 41705 14977 41739 15011
rect 42717 14977 42751 15011
rect 46029 14977 46063 15011
rect 47593 14977 47627 15011
rect 47869 14977 47903 15011
rect 51365 14977 51399 15011
rect 51549 14977 51583 15011
rect 52929 14977 52963 15011
rect 53205 14977 53239 15011
rect 54309 14977 54343 15011
rect 7389 14909 7423 14943
rect 10977 14909 11011 14943
rect 11621 14909 11655 14943
rect 12173 14909 12207 14943
rect 12449 14909 12483 14943
rect 17509 14909 17543 14943
rect 18981 14909 19015 14943
rect 19257 14909 19291 14943
rect 29009 14909 29043 14943
rect 30757 14909 30791 14943
rect 33885 14909 33919 14943
rect 40693 14909 40727 14943
rect 44833 14909 44867 14943
rect 45109 14909 45143 14943
rect 45293 14909 45327 14943
rect 45937 14909 45971 14943
rect 46857 14909 46891 14943
rect 47777 14909 47811 14943
rect 48973 14909 49007 14943
rect 51457 14909 51491 14943
rect 51641 14909 51675 14943
rect 53021 14909 53055 14943
rect 54217 14909 54251 14943
rect 56609 14909 56643 14943
rect 56885 14909 56919 14943
rect 9229 14841 9263 14875
rect 23121 14841 23155 14875
rect 54677 14841 54711 14875
rect 6745 14773 6779 14807
rect 8033 14773 8067 14807
rect 13921 14773 13955 14807
rect 24225 14773 24259 14807
rect 25973 14773 26007 14807
rect 28089 14773 28123 14807
rect 32229 14773 32263 14807
rect 36645 14773 36679 14807
rect 37289 14773 37323 14807
rect 41889 14773 41923 14807
rect 47593 14773 47627 14807
rect 48053 14773 48087 14807
rect 51181 14773 51215 14807
rect 53205 14773 53239 14807
rect 5917 14569 5951 14603
rect 6561 14569 6595 14603
rect 7665 14569 7699 14603
rect 9873 14569 9907 14603
rect 11909 14569 11943 14603
rect 13461 14569 13495 14603
rect 19625 14569 19659 14603
rect 29009 14569 29043 14603
rect 33885 14569 33919 14603
rect 46121 14569 46155 14603
rect 48513 14569 48547 14603
rect 53481 14569 53515 14603
rect 54125 14569 54159 14603
rect 58173 14569 58207 14603
rect 8309 14501 8343 14535
rect 12909 14501 12943 14535
rect 20361 14501 20395 14535
rect 26157 14501 26191 14535
rect 32873 14501 32907 14535
rect 43821 14501 43855 14535
rect 44373 14501 44407 14535
rect 45385 14501 45419 14535
rect 49065 14501 49099 14535
rect 51089 14501 51123 14535
rect 14289 14433 14323 14467
rect 21189 14433 21223 14467
rect 24409 14433 24443 14467
rect 24685 14433 24719 14467
rect 30573 14433 30607 14467
rect 36645 14433 36679 14467
rect 36921 14433 36955 14467
rect 39129 14433 39163 14467
rect 42625 14433 42659 14467
rect 45017 14433 45051 14467
rect 46213 14433 46247 14467
rect 46765 14433 46799 14467
rect 51825 14433 51859 14467
rect 53573 14433 53607 14467
rect 54309 14433 54343 14467
rect 56701 14433 56735 14467
rect 6653 14365 6687 14399
rect 7573 14365 7607 14399
rect 8217 14365 8251 14399
rect 9321 14365 9355 14399
rect 9781 14365 9815 14399
rect 12173 14365 12207 14399
rect 12725 14365 12759 14399
rect 13369 14365 13403 14399
rect 16037 14365 16071 14399
rect 16497 14365 16531 14399
rect 19533 14365 19567 14399
rect 20453 14365 20487 14399
rect 21097 14365 21131 14399
rect 22109 14365 22143 14399
rect 26801 14365 26835 14399
rect 27445 14365 27479 14399
rect 27629 14365 27663 14399
rect 29837 14365 29871 14399
rect 38117 14365 38151 14399
rect 38301 14365 38335 14399
rect 40325 14365 40359 14399
rect 40969 14365 41003 14399
rect 41245 14365 41279 14399
rect 41889 14365 41923 14399
rect 42901 14365 42935 14399
rect 43545 14365 43579 14399
rect 44465 14365 44499 14399
rect 45937 14365 45971 14399
rect 46029 14365 46063 14399
rect 46857 14365 46891 14399
rect 48237 14365 48271 14399
rect 48329 14365 48363 14399
rect 48973 14365 49007 14399
rect 49157 14365 49191 14399
rect 50721 14365 50755 14399
rect 51733 14365 51767 14399
rect 53297 14365 53331 14399
rect 53389 14365 53423 14399
rect 54033 14365 54067 14399
rect 56425 14365 56459 14399
rect 9229 14297 9263 14331
rect 15761 14297 15795 14331
rect 22385 14297 22419 14331
rect 30113 14297 30147 14331
rect 30849 14297 30883 14331
rect 48513 14297 48547 14331
rect 52561 14297 52595 14331
rect 52745 14297 52779 14331
rect 10425 14229 10459 14263
rect 17785 14229 17819 14263
rect 21465 14229 21499 14263
rect 23857 14229 23891 14263
rect 26709 14229 26743 14263
rect 28457 14229 28491 14263
rect 32321 14229 32355 14263
rect 35173 14229 35207 14263
rect 37565 14229 37599 14263
rect 40417 14229 40451 14263
rect 42165 14229 42199 14263
rect 45477 14229 45511 14263
rect 47225 14229 47259 14263
rect 48053 14229 48087 14263
rect 50537 14229 50571 14263
rect 50813 14229 50847 14263
rect 50905 14229 50939 14263
rect 52101 14229 52135 14263
rect 54309 14229 54343 14263
rect 6837 14025 6871 14059
rect 12265 14025 12299 14059
rect 12909 14025 12943 14059
rect 16129 14025 16163 14059
rect 17325 14025 17359 14059
rect 18521 14025 18555 14059
rect 23949 14025 23983 14059
rect 29561 14025 29595 14059
rect 33241 14025 33275 14059
rect 43637 14025 43671 14059
rect 45017 14025 45051 14059
rect 46121 14025 46155 14059
rect 46673 14025 46707 14059
rect 49341 14025 49375 14059
rect 50629 14025 50663 14059
rect 53849 14025 53883 14059
rect 54677 14025 54711 14059
rect 57253 14025 57287 14059
rect 21189 13957 21223 13991
rect 22477 13957 22511 13991
rect 30573 13957 30607 13991
rect 37749 13957 37783 13991
rect 44833 13957 44867 13991
rect 45109 13957 45143 13991
rect 47869 13957 47903 13991
rect 49801 13957 49835 13991
rect 49985 13957 50019 13991
rect 6745 13889 6779 13923
rect 7941 13889 7975 13923
rect 8769 13889 8803 13923
rect 11805 13889 11839 13923
rect 12449 13889 12483 13923
rect 13093 13889 13127 13923
rect 13829 13889 13863 13923
rect 16681 13889 16715 13923
rect 17417 13889 17451 13923
rect 18061 13889 18095 13923
rect 20269 13889 20303 13923
rect 21097 13889 21131 13923
rect 26985 13889 27019 13923
rect 27813 13889 27847 13923
rect 30297 13889 30331 13923
rect 31217 13889 31251 13923
rect 32413 13889 32447 13923
rect 33885 13889 33919 13923
rect 40049 13889 40083 13923
rect 40969 13889 41003 13923
rect 41705 13889 41739 13923
rect 42441 13889 42475 13923
rect 42717 13889 42751 13923
rect 43361 13889 43395 13923
rect 44281 13889 44315 13923
rect 45201 13889 45235 13923
rect 45385 13889 45419 13923
rect 45845 13889 45879 13923
rect 46581 13889 46615 13923
rect 46765 13889 46799 13923
rect 50537 13889 50571 13923
rect 50721 13889 50755 13923
rect 53205 13889 53239 13923
rect 53849 13889 53883 13923
rect 54033 13889 54067 13923
rect 54493 13889 54527 13923
rect 56241 13889 56275 13923
rect 58081 13889 58115 13923
rect 8033 13821 8067 13855
rect 9229 13821 9263 13855
rect 10977 13821 11011 13855
rect 11713 13821 11747 13855
rect 14381 13821 14415 13855
rect 22201 13821 22235 13855
rect 24409 13821 24443 13855
rect 26157 13821 26191 13855
rect 27077 13821 27111 13855
rect 28089 13821 28123 13855
rect 30573 13821 30607 13855
rect 31125 13821 31159 13855
rect 32689 13821 32723 13855
rect 34161 13821 34195 13855
rect 35633 13821 35667 13855
rect 37565 13821 37599 13855
rect 39405 13821 39439 13855
rect 40693 13821 40727 13855
rect 46121 13821 46155 13855
rect 47593 13821 47627 13855
rect 51365 13821 51399 13855
rect 51641 13821 51675 13855
rect 53389 13821 53423 13855
rect 56149 13821 56183 13855
rect 13645 13753 13679 13787
rect 17969 13753 18003 13787
rect 31585 13753 31619 13787
rect 40233 13753 40267 13787
rect 44097 13753 44131 13787
rect 45937 13753 45971 13787
rect 10713 13685 10747 13719
rect 14644 13685 14678 13719
rect 20005 13685 20039 13719
rect 24672 13685 24706 13719
rect 30389 13685 30423 13719
rect 41889 13685 41923 13719
rect 56517 13685 56551 13719
rect 57897 13685 57931 13719
rect 10057 13481 10091 13515
rect 12265 13481 12299 13515
rect 20361 13481 20395 13515
rect 24501 13481 24535 13515
rect 27353 13481 27387 13515
rect 28733 13481 28767 13515
rect 29653 13481 29687 13515
rect 33977 13481 34011 13515
rect 39313 13481 39347 13515
rect 40325 13481 40359 13515
rect 43821 13481 43855 13515
rect 46121 13481 46155 13515
rect 53389 13481 53423 13515
rect 58173 13481 58207 13515
rect 7205 13413 7239 13447
rect 19349 13413 19383 13447
rect 49157 13413 49191 13447
rect 7665 13345 7699 13379
rect 23857 13345 23891 13379
rect 30573 13345 30607 13379
rect 32689 13345 32723 13379
rect 37105 13345 37139 13379
rect 40969 13345 41003 13379
rect 42625 13345 42659 13379
rect 45293 13345 45327 13379
rect 45385 13345 45419 13379
rect 50261 13345 50295 13379
rect 51917 13345 51951 13379
rect 54217 13345 54251 13379
rect 56701 13345 56735 13379
rect 7573 13277 7607 13311
rect 11345 13277 11379 13311
rect 13553 13277 13587 13311
rect 16037 13277 16071 13311
rect 16865 13277 16899 13311
rect 19257 13277 19291 13311
rect 22109 13277 22143 13311
rect 24409 13277 24443 13311
rect 25605 13277 25639 13311
rect 28917 13277 28951 13311
rect 29745 13277 29779 13311
rect 30297 13277 30331 13311
rect 30389 13277 30423 13311
rect 32873 13277 32907 13311
rect 35679 13277 35713 13311
rect 37473 13277 37507 13311
rect 37933 13277 37967 13311
rect 40509 13277 40543 13311
rect 41245 13277 41279 13311
rect 41889 13277 41923 13311
rect 42901 13277 42935 13311
rect 43545 13277 43579 13311
rect 44281 13277 44315 13311
rect 44465 13277 44499 13311
rect 45477 13277 45511 13311
rect 45569 13277 45603 13311
rect 46305 13277 46339 13311
rect 47225 13277 47259 13311
rect 47409 13277 47443 13311
rect 47501 13277 47535 13311
rect 48237 13277 48271 13311
rect 50169 13277 50203 13311
rect 50353 13277 50387 13311
rect 50813 13277 50847 13311
rect 51641 13277 51675 13311
rect 54309 13277 54343 13311
rect 56425 13277 56459 13311
rect 15761 13209 15795 13243
rect 17049 13209 17083 13243
rect 18705 13209 18739 13243
rect 21649 13209 21683 13243
rect 26065 13209 26099 13243
rect 31033 13209 31067 13243
rect 34897 13209 34931 13243
rect 35081 13209 35115 13243
rect 42165 13209 42199 13243
rect 44373 13209 44407 13243
rect 48789 13209 48823 13243
rect 8309 13141 8343 13175
rect 9045 13141 9079 13175
rect 14289 13141 14323 13175
rect 25513 13141 25547 13175
rect 30573 13141 30607 13175
rect 33333 13141 33367 13175
rect 38117 13141 38151 13175
rect 45109 13141 45143 13175
rect 47041 13141 47075 13175
rect 48145 13141 48179 13175
rect 49249 13141 49283 13175
rect 50997 13141 51031 13175
rect 54677 13141 54711 13175
rect 9689 12937 9723 12971
rect 20913 12937 20947 12971
rect 25789 12937 25823 12971
rect 26985 12937 27019 12971
rect 30849 12937 30883 12971
rect 31017 12937 31051 12971
rect 35541 12937 35575 12971
rect 42625 12937 42659 12971
rect 50353 12937 50387 12971
rect 53389 12937 53423 12971
rect 53849 12937 53883 12971
rect 57345 12937 57379 12971
rect 58081 12937 58115 12971
rect 10977 12869 11011 12903
rect 14381 12869 14415 12903
rect 17325 12869 17359 12903
rect 22385 12869 22419 12903
rect 24501 12869 24535 12903
rect 29837 12869 29871 12903
rect 31217 12869 31251 12903
rect 51825 12869 51859 12903
rect 55321 12869 55355 12903
rect 7665 12801 7699 12835
rect 11805 12801 11839 12835
rect 12081 12801 12115 12835
rect 12633 12801 12667 12835
rect 13553 12801 13587 12835
rect 19901 12801 19935 12835
rect 20269 12801 20303 12835
rect 22109 12801 22143 12835
rect 27721 12801 27755 12835
rect 32321 12801 32355 12835
rect 33793 12801 33827 12835
rect 36001 12801 36035 12835
rect 37289 12801 37323 12835
rect 39129 12801 39163 12835
rect 40693 12801 40727 12835
rect 40969 12801 41003 12835
rect 41705 12801 41739 12835
rect 42441 12801 42475 12835
rect 44281 12801 44315 12835
rect 44741 12801 44775 12835
rect 44925 12801 44959 12835
rect 45477 12801 45511 12835
rect 46857 12801 46891 12835
rect 48329 12801 48363 12835
rect 49341 12801 49375 12835
rect 49433 12801 49467 12835
rect 53113 12801 53147 12835
rect 55597 12801 55631 12835
rect 56149 12801 56183 12835
rect 57161 12801 57195 12835
rect 57897 12801 57931 12835
rect 7757 12733 7791 12767
rect 13645 12733 13679 12767
rect 16129 12733 16163 12767
rect 17141 12733 17175 12767
rect 18613 12733 18647 12767
rect 28181 12733 28215 12767
rect 30021 12733 30055 12767
rect 32229 12733 32263 12767
rect 33149 12733 33183 12767
rect 34069 12733 34103 12767
rect 36093 12733 36127 12767
rect 37473 12733 37507 12767
rect 40141 12733 40175 12767
rect 41889 12733 41923 12767
rect 45661 12733 45695 12767
rect 48421 12733 48455 12767
rect 49157 12733 49191 12767
rect 52101 12733 52135 12767
rect 53389 12733 53423 12767
rect 13921 12665 13955 12699
rect 32689 12665 32723 12699
rect 46397 12665 46431 12699
rect 47041 12665 47075 12699
rect 48697 12665 48731 12699
rect 49249 12665 49283 12699
rect 53205 12665 53239 12699
rect 56333 12665 56367 12699
rect 7941 12597 7975 12631
rect 23857 12597 23891 12631
rect 27629 12597 27663 12631
rect 31033 12597 31067 12631
rect 36001 12597 36035 12631
rect 36369 12597 36403 12631
rect 39681 12597 39715 12631
rect 44833 12597 44867 12631
rect 47593 12597 47627 12631
rect 10885 12393 10919 12427
rect 14197 12393 14231 12427
rect 15117 12393 15151 12427
rect 23765 12393 23799 12427
rect 24409 12393 24443 12427
rect 30481 12393 30515 12427
rect 31033 12393 31067 12427
rect 39313 12393 39347 12427
rect 42165 12393 42199 12427
rect 46765 12393 46799 12427
rect 47225 12393 47259 12427
rect 51825 12393 51859 12427
rect 53113 12393 53147 12427
rect 53297 12393 53331 12427
rect 54125 12393 54159 12427
rect 54401 12393 54435 12427
rect 21281 12325 21315 12359
rect 28733 12325 28767 12359
rect 30297 12325 30331 12359
rect 34069 12325 34103 12359
rect 37197 12325 37231 12359
rect 49525 12325 49559 12359
rect 13277 12257 13311 12291
rect 25881 12257 25915 12291
rect 28457 12257 28491 12291
rect 32229 12257 32263 12291
rect 33609 12257 33643 12291
rect 34805 12257 34839 12291
rect 35449 12257 35483 12291
rect 37657 12257 37691 12291
rect 38209 12257 38243 12291
rect 40969 12257 41003 12291
rect 44005 12257 44039 12291
rect 48697 12257 48731 12291
rect 48973 12257 49007 12291
rect 52009 12257 52043 12291
rect 54033 12257 54067 12291
rect 57069 12257 57103 12291
rect 13185 12189 13219 12223
rect 16865 12189 16899 12223
rect 18705 12189 18739 12223
rect 19349 12189 19383 12223
rect 19717 12189 19751 12223
rect 23029 12189 23063 12223
rect 23857 12189 23891 12223
rect 26157 12189 26191 12223
rect 26709 12189 26743 12223
rect 26893 12189 26927 12223
rect 28365 12189 28399 12223
rect 30021 12189 30055 12223
rect 31217 12189 31251 12223
rect 31309 12189 31343 12223
rect 31953 12189 31987 12223
rect 33701 12189 33735 12223
rect 34713 12189 34747 12223
rect 34897 12189 34931 12223
rect 35725 12189 35759 12223
rect 37565 12189 37599 12223
rect 38393 12189 38427 12223
rect 38485 12189 38519 12223
rect 38669 12189 38703 12223
rect 38761 12189 38795 12223
rect 39865 12189 39899 12223
rect 40141 12189 40175 12223
rect 41245 12189 41279 12223
rect 41981 12189 42015 12223
rect 44097 12189 44131 12223
rect 45017 12189 45051 12223
rect 49433 12189 49467 12223
rect 49617 12189 49651 12223
rect 50445 12189 50479 12223
rect 50721 12189 50755 12223
rect 52101 12189 52135 12223
rect 54217 12189 54251 12223
rect 12173 12121 12207 12155
rect 16405 12121 16439 12155
rect 17049 12121 17083 12155
rect 22569 12121 22603 12155
rect 31033 12121 31067 12155
rect 42717 12121 42751 12155
rect 45293 12121 45327 12155
rect 53481 12121 53515 12155
rect 53941 12121 53975 12155
rect 56793 12121 56827 12155
rect 13553 12053 13587 12087
rect 20361 12053 20395 12087
rect 23121 12053 23155 12087
rect 27721 12053 27755 12087
rect 31493 12053 31527 12087
rect 39957 12053 39991 12087
rect 40325 12053 40359 12087
rect 42809 12053 42843 12087
rect 44465 12053 44499 12087
rect 53271 12053 53305 12087
rect 55321 12053 55355 12087
rect 12265 11849 12299 11883
rect 13277 11849 13311 11883
rect 14841 11849 14875 11883
rect 17877 11849 17911 11883
rect 18705 11849 18739 11883
rect 19625 11849 19659 11883
rect 25697 11849 25731 11883
rect 26249 11849 26283 11883
rect 30665 11849 30699 11883
rect 31493 11849 31527 11883
rect 33425 11849 33459 11883
rect 33793 11849 33827 11883
rect 35541 11849 35575 11883
rect 35725 11849 35759 11883
rect 40785 11849 40819 11883
rect 42625 11849 42659 11883
rect 53941 11849 53975 11883
rect 56609 11849 56643 11883
rect 13829 11781 13863 11815
rect 16129 11781 16163 11815
rect 16957 11781 16991 11815
rect 23765 11781 23799 11815
rect 28273 11781 28307 11815
rect 30757 11781 30791 11815
rect 43637 11781 43671 11815
rect 47961 11781 47995 11815
rect 54217 11781 54251 11815
rect 12633 11713 12667 11747
rect 18613 11713 18647 11747
rect 19717 11713 19751 11747
rect 20269 11713 20303 11747
rect 20637 11713 20671 11747
rect 22017 11713 22051 11747
rect 22201 11713 22235 11747
rect 23489 11713 23523 11747
rect 30573 11713 30607 11747
rect 31401 11713 31435 11747
rect 31585 11713 31619 11747
rect 32413 11713 32447 11747
rect 32597 11713 32631 11747
rect 33609 11713 33643 11747
rect 33885 11713 33919 11747
rect 34529 11713 34563 11747
rect 35357 11713 35391 11747
rect 35449 11713 35483 11747
rect 35725 11713 35759 11747
rect 36461 11713 36495 11747
rect 39957 11713 39991 11747
rect 40601 11713 40635 11747
rect 40785 11713 40819 11747
rect 41429 11713 41463 11747
rect 42441 11713 42475 11747
rect 44465 11713 44499 11747
rect 48145 11713 48179 11747
rect 48789 11713 48823 11747
rect 48973 11713 49007 11747
rect 50169 11713 50203 11747
rect 53113 11713 53147 11747
rect 53941 11713 53975 11747
rect 54033 11713 54067 11747
rect 54953 11713 54987 11747
rect 56241 11713 56275 11747
rect 12725 11645 12759 11679
rect 17417 11645 17451 11679
rect 21281 11645 21315 11679
rect 23029 11645 23063 11679
rect 28089 11645 28123 11679
rect 29929 11645 29963 11679
rect 30389 11645 30423 11679
rect 34437 11645 34471 11679
rect 37381 11645 37415 11679
rect 38853 11645 38887 11679
rect 39129 11645 39163 11679
rect 39589 11645 39623 11679
rect 39865 11645 39899 11679
rect 41337 11645 41371 11679
rect 44741 11645 44775 11679
rect 50813 11645 50847 11679
rect 51089 11645 51123 11679
rect 52929 11645 52963 11679
rect 53021 11645 53055 11679
rect 54861 11645 54895 11679
rect 56149 11645 56183 11679
rect 17693 11577 17727 11611
rect 30941 11577 30975 11611
rect 25237 11509 25271 11543
rect 32505 11509 32539 11543
rect 34805 11509 34839 11543
rect 36277 11509 36311 11543
rect 41705 11509 41739 11543
rect 43729 11509 43763 11543
rect 46213 11509 46247 11543
rect 48329 11509 48363 11543
rect 49157 11509 49191 11543
rect 50261 11509 50295 11543
rect 52101 11509 52135 11543
rect 53481 11509 53515 11543
rect 55229 11509 55263 11543
rect 12817 11305 12851 11339
rect 13553 11305 13587 11339
rect 14105 11305 14139 11339
rect 18429 11305 18463 11339
rect 24501 11305 24535 11339
rect 26985 11305 27019 11339
rect 28641 11305 28675 11339
rect 31585 11305 31619 11339
rect 32965 11305 32999 11339
rect 36829 11305 36863 11339
rect 38669 11305 38703 11339
rect 40417 11305 40451 11339
rect 45109 11305 45143 11339
rect 53205 11305 53239 11339
rect 56425 11305 56459 11339
rect 12265 11237 12299 11271
rect 40969 11237 41003 11271
rect 49433 11237 49467 11271
rect 52469 11237 52503 11271
rect 52561 11237 52595 11271
rect 53849 11237 53883 11271
rect 19349 11169 19383 11203
rect 19901 11169 19935 11203
rect 20177 11169 20211 11203
rect 22109 11169 22143 11203
rect 23857 11169 23891 11203
rect 29561 11169 29595 11203
rect 30021 11169 30055 11203
rect 30849 11169 30883 11203
rect 35357 11169 35391 11203
rect 37289 11169 37323 11203
rect 39037 11169 39071 11203
rect 40233 11169 40267 11203
rect 42717 11169 42751 11203
rect 45293 11169 45327 11203
rect 48329 11169 48363 11203
rect 48973 11169 49007 11203
rect 50445 11169 50479 11203
rect 52377 11169 52411 11203
rect 57897 11169 57931 11203
rect 58173 11169 58207 11203
rect 12173 11101 12207 11135
rect 15117 11101 15151 11135
rect 15761 11101 15795 11135
rect 18521 11101 18555 11135
rect 19441 11101 19475 11135
rect 24593 11101 24627 11135
rect 25421 11101 25455 11135
rect 25605 11101 25639 11135
rect 28549 11101 28583 11135
rect 28733 11101 28767 11135
rect 29745 11101 29779 11135
rect 29837 11101 29871 11135
rect 29929 11101 29963 11135
rect 30757 11101 30791 11135
rect 30941 11101 30975 11135
rect 32505 11101 32539 11135
rect 32597 11101 32631 11135
rect 32781 11101 32815 11135
rect 35081 11101 35115 11135
rect 38117 11101 38151 11135
rect 38945 11101 38979 11135
rect 40141 11101 40175 11135
rect 45385 11101 45419 11135
rect 47225 11101 47259 11135
rect 47409 11101 47443 11135
rect 47869 11101 47903 11135
rect 48145 11101 48179 11135
rect 49065 11101 49099 11135
rect 50169 11101 50203 11135
rect 52653 11101 52687 11135
rect 53113 11101 53147 11135
rect 53297 11101 53331 11135
rect 53941 11101 53975 11135
rect 16037 11033 16071 11067
rect 22385 11033 22419 11067
rect 28089 11033 28123 11067
rect 31493 11033 31527 11067
rect 33517 11033 33551 11067
rect 34069 11033 34103 11067
rect 42441 11033 42475 11067
rect 47317 11033 47351 11067
rect 47961 11033 47995 11067
rect 15209 10965 15243 10999
rect 17509 10965 17543 10999
rect 21649 10965 21683 10999
rect 26433 10965 26467 10999
rect 43545 10965 43579 10999
rect 51917 10965 51951 10999
rect 1961 10761 1995 10795
rect 16129 10761 16163 10795
rect 17141 10761 17175 10795
rect 21189 10761 21223 10795
rect 26433 10761 26467 10795
rect 36369 10761 36403 10795
rect 42441 10761 42475 10795
rect 43269 10761 43303 10795
rect 48881 10761 48915 10795
rect 49433 10761 49467 10795
rect 52009 10761 52043 10795
rect 17693 10693 17727 10727
rect 20453 10693 20487 10727
rect 22201 10693 22235 10727
rect 24593 10693 24627 10727
rect 29745 10693 29779 10727
rect 33793 10693 33827 10727
rect 35541 10693 35575 10727
rect 39037 10693 39071 10727
rect 41245 10693 41279 10727
rect 41429 10693 41463 10727
rect 49709 10693 49743 10727
rect 51733 10693 51767 10727
rect 1869 10625 1903 10659
rect 20729 10625 20763 10659
rect 21925 10625 21959 10659
rect 25421 10625 25455 10659
rect 25605 10625 25639 10659
rect 32321 10625 32355 10659
rect 36553 10625 36587 10659
rect 37749 10625 37783 10659
rect 37841 10625 37875 10659
rect 38393 10625 38427 10659
rect 42717 10625 42751 10659
rect 43361 10625 43395 10659
rect 44281 10625 44315 10659
rect 48697 10625 48731 10659
rect 48973 10625 49007 10659
rect 49433 10625 49467 10659
rect 49525 10625 49559 10659
rect 51641 10625 51675 10659
rect 51825 10625 51859 10659
rect 53021 10625 53055 10659
rect 14381 10557 14415 10591
rect 14657 10557 14691 10591
rect 16681 10557 16715 10591
rect 18981 10557 19015 10591
rect 24317 10557 24351 10591
rect 24777 10557 24811 10591
rect 27169 10557 27203 10591
rect 28641 10557 28675 10591
rect 28825 10557 28859 10591
rect 29561 10557 29595 10591
rect 30757 10557 30791 10591
rect 32229 10557 32263 10591
rect 37565 10557 37599 10591
rect 38577 10557 38611 10591
rect 42441 10557 42475 10591
rect 44005 10557 44039 10591
rect 52929 10557 52963 10591
rect 17049 10489 17083 10523
rect 42625 10489 42659 10523
rect 48513 10489 48547 10523
rect 51457 10489 51491 10523
rect 53389 10489 53423 10523
rect 13829 10421 13863 10455
rect 18521 10421 18555 10455
rect 32597 10421 32631 10455
rect 37841 10421 37875 10455
rect 40325 10421 40359 10455
rect 45385 10421 45419 10455
rect 47685 10421 47719 10455
rect 1593 10217 1627 10251
rect 16221 10217 16255 10251
rect 19625 10217 19659 10251
rect 30665 10217 30699 10251
rect 31217 10217 31251 10251
rect 31493 10217 31527 10251
rect 34970 10217 35004 10251
rect 40601 10217 40635 10251
rect 45569 10217 45603 10251
rect 48329 10217 48363 10251
rect 52377 10217 52411 10251
rect 52837 10217 52871 10251
rect 21097 10149 21131 10183
rect 29837 10149 29871 10183
rect 33241 10149 33275 10183
rect 55873 10149 55907 10183
rect 18153 10081 18187 10115
rect 23857 10081 23891 10115
rect 26525 10081 26559 10115
rect 26709 10081 26743 10115
rect 27169 10081 27203 10115
rect 28825 10081 28859 10115
rect 29009 10081 29043 10115
rect 30021 10081 30055 10115
rect 30573 10081 30607 10115
rect 30757 10081 30791 10115
rect 31493 10081 31527 10115
rect 34713 10081 34747 10115
rect 36921 10081 36955 10115
rect 38669 10081 38703 10115
rect 40049 10081 40083 10115
rect 43269 10081 43303 10115
rect 51089 10081 51123 10115
rect 52469 10081 52503 10115
rect 56333 10081 56367 10115
rect 58081 10081 58115 10115
rect 19533 10013 19567 10047
rect 21189 10013 21223 10047
rect 22109 10013 22143 10047
rect 30481 10013 30515 10047
rect 31408 10013 31442 10047
rect 32689 10013 32723 10047
rect 39129 10013 39163 10047
rect 39313 10013 39347 10047
rect 51365 10013 51399 10047
rect 52377 10013 52411 10047
rect 52653 10013 52687 10047
rect 20361 9945 20395 9979
rect 24869 9945 24903 9979
rect 29561 9945 29595 9979
rect 31677 9945 31711 9979
rect 32229 9945 32263 9979
rect 34069 9945 34103 9979
rect 37197 9945 37231 9979
rect 39221 9945 39255 9979
rect 42993 9945 43027 9979
rect 45477 9945 45511 9979
rect 57805 9945 57839 9979
rect 15577 9877 15611 9911
rect 17509 9877 17543 9911
rect 18705 9877 18739 9911
rect 20269 9877 20303 9911
rect 33977 9877 34011 9911
rect 36461 9877 36495 9911
rect 40141 9877 40175 9911
rect 40233 9877 40267 9911
rect 41521 9877 41555 9911
rect 43821 9877 43855 9911
rect 44281 9877 44315 9911
rect 40759 9673 40793 9707
rect 43545 9673 43579 9707
rect 20729 9605 20763 9639
rect 21833 9605 21867 9639
rect 25881 9605 25915 9639
rect 28641 9605 28675 9639
rect 29929 9605 29963 9639
rect 38393 9605 38427 9639
rect 40969 9605 41003 9639
rect 41613 9605 41647 9639
rect 51825 9605 51859 9639
rect 52009 9605 52043 9639
rect 54585 9605 54619 9639
rect 58081 9605 58115 9639
rect 20821 9537 20855 9571
rect 32689 9537 32723 9571
rect 33701 9537 33735 9571
rect 36185 9537 36219 9571
rect 37473 9537 37507 9571
rect 42625 9537 42659 9571
rect 44465 9537 44499 9571
rect 47777 9537 47811 9571
rect 48881 9537 48915 9571
rect 54309 9537 54343 9571
rect 18429 9469 18463 9503
rect 18705 9469 18739 9503
rect 24685 9469 24719 9503
rect 26065 9469 26099 9503
rect 27445 9469 27479 9503
rect 28825 9469 28859 9503
rect 29745 9469 29779 9503
rect 30665 9469 30699 9503
rect 33977 9469 34011 9503
rect 37289 9469 37323 9503
rect 42533 9469 42567 9503
rect 47869 9469 47903 9503
rect 49157 9469 49191 9503
rect 50629 9469 50663 9503
rect 56057 9469 56091 9503
rect 32505 9401 32539 9435
rect 36001 9401 36035 9435
rect 40601 9401 40635 9435
rect 44649 9401 44683 9435
rect 48145 9401 48179 9435
rect 17877 9333 17911 9367
rect 20177 9333 20211 9367
rect 35449 9333 35483 9367
rect 39681 9333 39715 9367
rect 40785 9333 40819 9367
rect 41521 9333 41555 9367
rect 42901 9333 42935 9367
rect 3249 9129 3283 9163
rect 18613 9129 18647 9163
rect 19533 9129 19567 9163
rect 21005 9129 21039 9163
rect 26709 9129 26743 9163
rect 35173 9129 35207 9163
rect 40325 9129 40359 9163
rect 41245 9129 41279 9163
rect 42735 9129 42769 9163
rect 48237 9129 48271 9163
rect 50353 9129 50387 9163
rect 20269 9061 20303 9095
rect 25789 9061 25823 9095
rect 30113 9061 30147 9095
rect 36829 9061 36863 9095
rect 43729 9061 43763 9095
rect 26525 8993 26559 9027
rect 27353 8993 27387 9027
rect 27905 8993 27939 9027
rect 28273 8993 28307 9027
rect 28365 8993 28399 9027
rect 29653 8993 29687 9027
rect 31033 8993 31067 9027
rect 31585 8993 31619 9027
rect 38117 8993 38151 9027
rect 38945 8993 38979 9027
rect 40233 8993 40267 9027
rect 42993 8993 43027 9027
rect 45661 8993 45695 9027
rect 57069 8993 57103 9027
rect 57345 8993 57379 9027
rect 2697 8925 2731 8959
rect 16865 8925 16899 8959
rect 26433 8925 26467 8959
rect 27261 8925 27295 8959
rect 27445 8925 27479 8959
rect 28089 8925 28123 8959
rect 28181 8925 28215 8959
rect 29745 8925 29779 8959
rect 31401 8925 31435 8959
rect 32413 8925 32447 8959
rect 35173 8925 35207 8959
rect 35265 8925 35299 8959
rect 36461 8925 36495 8959
rect 37841 8925 37875 8959
rect 38761 8925 38795 8959
rect 38853 8925 38887 8959
rect 39037 8925 39071 8959
rect 40049 8925 40083 8959
rect 40325 8925 40359 8959
rect 43545 8925 43579 8959
rect 45569 8925 45603 8959
rect 50169 8925 50203 8959
rect 17141 8857 17175 8891
rect 19993 8857 20027 8891
rect 29009 8857 29043 8891
rect 31309 8857 31343 8891
rect 32689 8857 32723 8891
rect 35449 8857 35483 8891
rect 36553 8857 36587 8891
rect 44373 8857 44407 8891
rect 50997 8857 51031 8891
rect 2513 8789 2547 8823
rect 16313 8789 16347 8823
rect 20453 8789 20487 8823
rect 21465 8789 21499 8823
rect 31217 8789 31251 8823
rect 34161 8789 34195 8823
rect 34989 8789 35023 8823
rect 36277 8789 36311 8823
rect 36645 8789 36679 8823
rect 38577 8789 38611 8823
rect 39865 8789 39899 8823
rect 44281 8789 44315 8823
rect 45201 8789 45235 8823
rect 46305 8789 46339 8823
rect 55597 8789 55631 8823
rect 18705 8585 18739 8619
rect 28825 8585 28859 8619
rect 29377 8585 29411 8619
rect 30389 8585 30423 8619
rect 31493 8585 31527 8619
rect 32689 8585 32723 8619
rect 33471 8585 33505 8619
rect 36369 8585 36403 8619
rect 40969 8585 41003 8619
rect 42441 8585 42475 8619
rect 45293 8585 45327 8619
rect 45477 8585 45511 8619
rect 46213 8585 46247 8619
rect 55413 8585 55447 8619
rect 19901 8517 19935 8551
rect 27353 8517 27387 8551
rect 27905 8517 27939 8551
rect 43177 8517 43211 8551
rect 45661 8517 45695 8551
rect 21005 8449 21039 8483
rect 28457 8449 28491 8483
rect 29285 8449 29319 8483
rect 29469 8449 29503 8483
rect 30573 8449 30607 8483
rect 30665 8449 30699 8483
rect 30849 8449 30883 8483
rect 30941 8449 30975 8483
rect 32321 8449 32355 8483
rect 35265 8449 35299 8483
rect 36277 8449 36311 8483
rect 36553 8449 36587 8483
rect 37473 8449 37507 8483
rect 38563 8449 38597 8483
rect 39865 8449 39899 8483
rect 40693 8449 40727 8483
rect 40785 8449 40819 8483
rect 41613 8449 41647 8483
rect 44373 8449 44407 8483
rect 44649 8449 44683 8483
rect 45385 8449 45419 8483
rect 46397 8449 46431 8483
rect 46581 8449 46615 8483
rect 46673 8449 46707 8483
rect 20361 8381 20395 8415
rect 28549 8381 28583 8415
rect 32229 8381 32263 8415
rect 34897 8381 34931 8415
rect 36737 8381 36771 8415
rect 37381 8381 37415 8415
rect 38393 8381 38427 8415
rect 39957 8381 39991 8415
rect 40969 8381 41003 8415
rect 44557 8381 44591 8415
rect 20177 8313 20211 8347
rect 20821 8313 20855 8347
rect 35817 8313 35851 8347
rect 37841 8313 37875 8347
rect 38853 8313 38887 8347
rect 41429 8313 41463 8347
rect 44189 8313 44223 8347
rect 45109 8313 45143 8347
rect 28457 8245 28491 8279
rect 40233 8245 40267 8279
rect 43085 8245 43119 8279
rect 44373 8245 44407 8279
rect 21189 8041 21223 8075
rect 26893 8041 26927 8075
rect 28089 8041 28123 8075
rect 30849 8041 30883 8075
rect 32781 8041 32815 8075
rect 37013 8041 37047 8075
rect 41889 8041 41923 8075
rect 47317 8041 47351 8075
rect 29837 7973 29871 8007
rect 31677 7973 31711 8007
rect 39313 7973 39347 8007
rect 45017 7973 45051 8007
rect 57897 7973 57931 8007
rect 27905 7905 27939 7939
rect 29009 7905 29043 7939
rect 30573 7905 30607 7939
rect 34713 7905 34747 7939
rect 36461 7905 36495 7939
rect 38485 7905 38519 7939
rect 38761 7905 38795 7939
rect 40141 7905 40175 7939
rect 42349 7905 42383 7939
rect 42625 7905 42659 7939
rect 45477 7905 45511 7939
rect 46029 7905 46063 7939
rect 20361 7837 20395 7871
rect 20545 7837 20579 7871
rect 28089 7837 28123 7871
rect 28733 7837 28767 7871
rect 28825 7837 28859 7871
rect 30481 7837 30515 7871
rect 32321 7837 32355 7871
rect 32597 7837 32631 7871
rect 33701 7837 33735 7871
rect 33977 7837 34011 7871
rect 45385 7837 45419 7871
rect 46213 7837 46247 7871
rect 46489 7837 46523 7871
rect 46949 7837 46983 7871
rect 27813 7769 27847 7803
rect 29009 7769 29043 7803
rect 31401 7769 31435 7803
rect 32413 7769 32447 7803
rect 34989 7769 35023 7803
rect 40417 7769 40451 7803
rect 47133 7769 47167 7803
rect 57437 7769 57471 7803
rect 58081 7769 58115 7803
rect 20729 7701 20763 7735
rect 28273 7701 28307 7735
rect 31861 7701 31895 7735
rect 33793 7701 33827 7735
rect 34161 7701 34195 7735
rect 44097 7701 44131 7735
rect 46397 7701 46431 7735
rect 27353 7497 27387 7531
rect 29009 7497 29043 7531
rect 29929 7497 29963 7531
rect 32689 7497 32723 7531
rect 37657 7497 37691 7531
rect 41337 7497 41371 7531
rect 44189 7497 44223 7531
rect 44741 7497 44775 7531
rect 46121 7497 46155 7531
rect 46581 7497 46615 7531
rect 22017 7429 22051 7463
rect 29177 7429 29211 7463
rect 29377 7429 29411 7463
rect 33517 7429 33551 7463
rect 33701 7429 33735 7463
rect 39773 7429 39807 7463
rect 40785 7429 40819 7463
rect 45753 7429 45787 7463
rect 46673 7429 46707 7463
rect 46857 7429 46891 7463
rect 20913 7361 20947 7395
rect 27537 7361 27571 7395
rect 28273 7361 28307 7395
rect 29837 7361 29871 7395
rect 30021 7361 30055 7395
rect 31125 7361 31159 7395
rect 32321 7361 32355 7395
rect 34437 7361 34471 7395
rect 37565 7361 37599 7395
rect 37749 7361 37783 7395
rect 40049 7361 40083 7395
rect 40601 7361 40635 7395
rect 41429 7361 41463 7395
rect 42441 7361 42475 7395
rect 44649 7361 44683 7395
rect 45937 7361 45971 7395
rect 46581 7361 46615 7395
rect 21925 7293 21959 7327
rect 28089 7293 28123 7327
rect 28181 7293 28215 7327
rect 28365 7293 28399 7327
rect 31217 7293 31251 7327
rect 32229 7293 32263 7327
rect 34345 7293 34379 7327
rect 38301 7293 38335 7327
rect 42717 7293 42751 7327
rect 21097 7225 21131 7259
rect 22477 7225 22511 7259
rect 31493 7225 31527 7259
rect 36737 7225 36771 7259
rect 28549 7157 28583 7191
rect 29193 7157 29227 7191
rect 34713 7157 34747 7191
rect 21649 6953 21683 6987
rect 30573 6953 30607 6987
rect 31585 6953 31619 6987
rect 31677 6953 31711 6987
rect 33517 6953 33551 6987
rect 35614 6953 35648 6987
rect 45109 6953 45143 6987
rect 45937 6953 45971 6987
rect 46489 6953 46523 6987
rect 27997 6885 28031 6919
rect 20361 6817 20395 6851
rect 31493 6817 31527 6851
rect 32229 6817 32263 6851
rect 37105 6817 37139 6851
rect 39037 6817 39071 6851
rect 40969 6817 41003 6851
rect 20177 6749 20211 6783
rect 27353 6749 27387 6783
rect 27537 6749 27571 6783
rect 28181 6749 28215 6783
rect 29561 6749 29595 6783
rect 29745 6749 29779 6783
rect 30481 6749 30515 6783
rect 30573 6749 30607 6783
rect 30849 6749 30883 6783
rect 31769 6749 31803 6783
rect 33425 6749 33459 6783
rect 33609 6749 33643 6783
rect 34713 6749 34747 6783
rect 35357 6749 35391 6783
rect 38209 6749 38243 6783
rect 38945 6749 38979 6783
rect 39129 6749 39163 6783
rect 40417 6749 40451 6783
rect 41797 6749 41831 6783
rect 41981 6749 42015 6783
rect 42625 6749 42659 6783
rect 45845 6749 45879 6783
rect 46029 6749 46063 6783
rect 47041 6749 47075 6783
rect 28365 6681 28399 6715
rect 38025 6681 38059 6715
rect 42441 6681 42475 6715
rect 43821 6681 43855 6715
rect 19717 6613 19751 6647
rect 27445 6613 27479 6647
rect 28273 6613 28307 6647
rect 28549 6613 28583 6647
rect 29745 6613 29779 6647
rect 30665 6613 30699 6647
rect 40325 6613 40359 6647
rect 41889 6613 41923 6647
rect 42809 6613 42843 6647
rect 43729 6613 43763 6647
rect 19533 6409 19567 6443
rect 35081 6409 35115 6443
rect 36737 6409 36771 6443
rect 42809 6409 42843 6443
rect 45661 6409 45695 6443
rect 46121 6409 46155 6443
rect 27169 6341 27203 6375
rect 28181 6341 28215 6375
rect 33609 6341 33643 6375
rect 41153 6341 41187 6375
rect 44649 6341 44683 6375
rect 27721 6273 27755 6307
rect 29377 6273 29411 6307
rect 31033 6273 31067 6307
rect 37749 6273 37783 6307
rect 37933 6273 37967 6307
rect 38761 6273 38795 6307
rect 39037 6273 39071 6307
rect 40233 6273 40267 6307
rect 41705 6273 41739 6307
rect 42717 6273 42751 6307
rect 42993 6273 43027 6307
rect 44005 6273 44039 6307
rect 27077 6205 27111 6239
rect 29101 6205 29135 6239
rect 30941 6205 30975 6239
rect 33333 6205 33367 6239
rect 38853 6205 38887 6239
rect 40325 6205 40359 6239
rect 40969 6205 41003 6239
rect 43177 6205 43211 6239
rect 43913 6205 43947 6239
rect 28457 6137 28491 6171
rect 28641 6137 28675 6171
rect 29285 6137 29319 6171
rect 31401 6137 31435 6171
rect 39221 6137 39255 6171
rect 43637 6137 43671 6171
rect 29193 6069 29227 6103
rect 29929 6069 29963 6103
rect 37841 6069 37875 6103
rect 39037 6069 39071 6103
rect 39865 6069 39899 6103
rect 41889 6069 41923 6103
rect 25973 5865 26007 5899
rect 27905 5865 27939 5899
rect 39865 5865 39899 5899
rect 29009 5797 29043 5831
rect 36369 5797 36403 5831
rect 39037 5797 39071 5831
rect 44097 5797 44131 5831
rect 28733 5729 28767 5763
rect 32413 5729 32447 5763
rect 32689 5729 32723 5763
rect 37289 5729 37323 5763
rect 40509 5729 40543 5763
rect 41337 5729 41371 5763
rect 42349 5729 42383 5763
rect 25789 5661 25823 5695
rect 28641 5661 28675 5695
rect 30481 5661 30515 5695
rect 30757 5661 30791 5695
rect 31401 5661 31435 5695
rect 40325 5661 40359 5695
rect 41245 5661 41279 5695
rect 42533 5661 42567 5695
rect 42717 5661 42751 5695
rect 42809 5661 42843 5695
rect 43637 5661 43671 5695
rect 44097 5661 44131 5695
rect 31217 5593 31251 5627
rect 35081 5593 35115 5627
rect 37565 5593 37599 5627
rect 43269 5593 43303 5627
rect 43453 5593 43487 5627
rect 44189 5593 44223 5627
rect 44373 5593 44407 5627
rect 30297 5525 30331 5559
rect 30665 5525 30699 5559
rect 34161 5525 34195 5559
rect 40233 5525 40267 5559
rect 41613 5525 41647 5559
rect 20637 5321 20671 5355
rect 21833 5321 21867 5355
rect 26249 5321 26283 5355
rect 30941 5321 30975 5355
rect 33333 5321 33367 5355
rect 37289 5321 37323 5355
rect 40325 5321 40359 5355
rect 41429 5321 41463 5355
rect 35725 5253 35759 5287
rect 39037 5253 39071 5287
rect 41613 5253 41647 5287
rect 41797 5253 41831 5287
rect 1685 5185 1719 5219
rect 21097 5185 21131 5219
rect 25881 5185 25915 5219
rect 26065 5185 26099 5219
rect 28733 5185 28767 5219
rect 29837 5185 29871 5219
rect 30849 5185 30883 5219
rect 31033 5185 31067 5219
rect 32321 5185 32355 5219
rect 32505 5185 32539 5219
rect 32597 5185 32631 5219
rect 37657 5185 37691 5219
rect 38577 5185 38611 5219
rect 41245 5185 41279 5219
rect 41521 5185 41555 5219
rect 42625 5185 42659 5219
rect 42901 5185 42935 5219
rect 21281 5117 21315 5151
rect 28825 5117 28859 5151
rect 29561 5117 29595 5151
rect 34805 5117 34839 5151
rect 35081 5117 35115 5151
rect 37749 5117 37783 5151
rect 38301 5117 38335 5151
rect 42717 5117 42751 5151
rect 2237 5049 2271 5083
rect 29101 5049 29135 5083
rect 35541 5049 35575 5083
rect 1501 4981 1535 5015
rect 25053 4981 25087 5015
rect 32137 4981 32171 5015
rect 38393 4981 38427 5015
rect 38485 4981 38519 5015
rect 42441 4981 42475 5015
rect 42901 4981 42935 5015
rect 24777 4777 24811 4811
rect 25881 4777 25915 4811
rect 31033 4777 31067 4811
rect 31953 4777 31987 4811
rect 33977 4777 34011 4811
rect 37565 4777 37599 4811
rect 39957 4777 39991 4811
rect 41705 4777 41739 4811
rect 25789 4709 25823 4743
rect 26617 4709 26651 4743
rect 33333 4709 33367 4743
rect 33425 4709 33459 4743
rect 38485 4709 38519 4743
rect 41153 4709 41187 4743
rect 27261 4641 27295 4675
rect 28733 4641 28767 4675
rect 30849 4641 30883 4675
rect 33241 4641 33275 4675
rect 38209 4641 38243 4675
rect 38393 4641 38427 4675
rect 43453 4641 43487 4675
rect 24869 4573 24903 4607
rect 29009 4573 29043 4607
rect 30757 4573 30791 4607
rect 31861 4573 31895 4607
rect 32045 4573 32079 4607
rect 33517 4573 33551 4607
rect 38485 4573 38519 4607
rect 40049 4573 40083 4607
rect 25421 4505 25455 4539
rect 26341 4505 26375 4539
rect 35081 4505 35115 4539
rect 35265 4505 35299 4539
rect 37549 4505 37583 4539
rect 37749 4505 37783 4539
rect 43177 4505 43211 4539
rect 26801 4437 26835 4471
rect 29653 4437 29687 4471
rect 37381 4437 37415 4471
rect 26985 4233 27019 4267
rect 40601 4233 40635 4267
rect 39129 4165 39163 4199
rect 27169 4097 27203 4131
rect 31033 4097 31067 4131
rect 32689 4097 32723 4131
rect 37473 4097 37507 4131
rect 42441 4097 42475 4131
rect 48697 4097 48731 4131
rect 49341 4097 49375 4131
rect 24593 4029 24627 4063
rect 24869 4029 24903 4063
rect 31125 4029 31159 4063
rect 32965 4029 32999 4063
rect 34897 4029 34931 4063
rect 35173 4029 35207 4063
rect 36645 4029 36679 4063
rect 37565 4029 37599 4063
rect 38853 4029 38887 4063
rect 42717 4029 42751 4063
rect 44189 4029 44223 4063
rect 31401 3961 31435 3995
rect 37841 3961 37875 3995
rect 23121 3893 23155 3927
rect 25329 3893 25363 3927
rect 29193 3893 29227 3927
rect 34437 3893 34471 3927
rect 48881 3893 48915 3927
rect 27169 3689 27203 3723
rect 27721 3689 27755 3723
rect 34713 3621 34747 3655
rect 41613 3621 41647 3655
rect 25697 3553 25731 3587
rect 36461 3553 36495 3587
rect 39865 3553 39899 3587
rect 25421 3485 25455 3519
rect 36185 3417 36219 3451
rect 40141 3417 40175 3451
rect 14197 3145 14231 3179
rect 37289 3145 37323 3179
rect 38761 3077 38795 3111
rect 19809 3009 19843 3043
rect 27905 3009 27939 3043
rect 28549 3009 28583 3043
rect 33333 3009 33367 3043
rect 57897 3009 57931 3043
rect 39037 2941 39071 2975
rect 39497 2941 39531 2975
rect 28089 2873 28123 2907
rect 19625 2805 19659 2839
rect 33517 2805 33551 2839
rect 52929 2805 52963 2839
rect 58081 2805 58115 2839
rect 38209 2601 38243 2635
rect 43269 2601 43303 2635
rect 10057 2533 10091 2567
rect 53113 2533 53147 2567
rect 1685 2397 1719 2431
rect 4169 2397 4203 2431
rect 4629 2397 4663 2431
rect 14289 2397 14323 2431
rect 19717 2397 19751 2431
rect 24685 2397 24719 2431
rect 29561 2397 29595 2431
rect 33793 2397 33827 2431
rect 38761 2397 38795 2431
rect 43453 2397 43487 2431
rect 43913 2397 43947 2431
rect 48421 2397 48455 2431
rect 57897 2397 57931 2431
rect 9321 2329 9355 2363
rect 9873 2329 9907 2363
rect 25237 2329 25271 2363
rect 53297 2329 53331 2363
rect 1501 2261 1535 2295
rect 4813 2261 4847 2295
rect 14473 2261 14507 2295
rect 19533 2261 19567 2295
rect 24501 2261 24535 2295
rect 29745 2261 29779 2295
rect 33609 2261 33643 2295
rect 38945 2261 38979 2295
rect 48605 2261 48639 2295
rect 58081 2261 58115 2295
<< metal1 >>
rect 1104 33754 58880 33776
rect 1104 33702 15398 33754
rect 15450 33702 15462 33754
rect 15514 33702 15526 33754
rect 15578 33702 15590 33754
rect 15642 33702 15654 33754
rect 15706 33702 29846 33754
rect 29898 33702 29910 33754
rect 29962 33702 29974 33754
rect 30026 33702 30038 33754
rect 30090 33702 30102 33754
rect 30154 33702 44294 33754
rect 44346 33702 44358 33754
rect 44410 33702 44422 33754
rect 44474 33702 44486 33754
rect 44538 33702 44550 33754
rect 44602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1486 33640 1492 33652
rect 1447 33612 1492 33640
rect 1486 33600 1492 33612
rect 1544 33600 1550 33652
rect 4798 33640 4804 33652
rect 4759 33612 4804 33640
rect 4798 33600 4804 33612
rect 4856 33600 4862 33652
rect 9030 33600 9036 33652
rect 9088 33640 9094 33652
rect 9217 33643 9275 33649
rect 9217 33640 9229 33643
rect 9088 33612 9229 33640
rect 9088 33600 9094 33612
rect 9217 33609 9229 33612
rect 9263 33609 9275 33643
rect 14366 33640 14372 33652
rect 14327 33612 14372 33640
rect 9217 33603 9275 33609
rect 14366 33600 14372 33612
rect 14424 33600 14430 33652
rect 18690 33600 18696 33652
rect 18748 33640 18754 33652
rect 19245 33643 19303 33649
rect 19245 33640 19257 33643
rect 18748 33612 19257 33640
rect 18748 33600 18754 33612
rect 19245 33609 19257 33612
rect 19291 33609 19303 33643
rect 33778 33640 33784 33652
rect 33739 33612 33784 33640
rect 19245 33603 19303 33609
rect 33778 33600 33784 33612
rect 33836 33600 33842 33652
rect 38654 33600 38660 33652
rect 38712 33640 38718 33652
rect 38749 33643 38807 33649
rect 38749 33640 38761 33643
rect 38712 33612 38761 33640
rect 38712 33600 38718 33612
rect 38749 33609 38761 33612
rect 38795 33609 38807 33643
rect 43254 33640 43260 33652
rect 43215 33612 43260 33640
rect 38749 33603 38807 33609
rect 43254 33600 43260 33612
rect 43312 33600 43318 33652
rect 48590 33640 48596 33652
rect 48551 33612 48596 33640
rect 48590 33600 48596 33612
rect 48648 33600 48654 33652
rect 53098 33640 53104 33652
rect 53059 33612 53104 33640
rect 53098 33600 53104 33612
rect 53156 33600 53162 33652
rect 27985 33575 28043 33581
rect 27985 33541 27997 33575
rect 28031 33572 28043 33575
rect 28534 33572 28540 33584
rect 28031 33544 28540 33572
rect 28031 33541 28043 33544
rect 27985 33535 28043 33541
rect 28534 33532 28540 33544
rect 28592 33532 28598 33584
rect 1670 33504 1676 33516
rect 1631 33476 1676 33504
rect 1670 33464 1676 33476
rect 1728 33464 1734 33516
rect 4614 33504 4620 33516
rect 4575 33476 4620 33504
rect 4614 33464 4620 33476
rect 4672 33464 4678 33516
rect 9398 33504 9404 33516
rect 9359 33476 9404 33504
rect 9398 33464 9404 33476
rect 9456 33464 9462 33516
rect 14553 33507 14611 33513
rect 14553 33473 14565 33507
rect 14599 33504 14611 33507
rect 17218 33504 17224 33516
rect 14599 33476 17224 33504
rect 14599 33473 14611 33476
rect 14553 33467 14611 33473
rect 17218 33464 17224 33476
rect 17276 33464 17282 33516
rect 19426 33504 19432 33516
rect 19387 33476 19432 33504
rect 19426 33464 19432 33476
rect 19484 33464 19490 33516
rect 23842 33464 23848 33516
rect 23900 33504 23906 33516
rect 24581 33507 24639 33513
rect 24581 33504 24593 33507
rect 23900 33476 24593 33504
rect 23900 33464 23906 33476
rect 24581 33473 24593 33476
rect 24627 33504 24639 33507
rect 25041 33507 25099 33513
rect 25041 33504 25053 33507
rect 24627 33476 25053 33504
rect 24627 33473 24639 33476
rect 24581 33467 24639 33473
rect 25041 33473 25053 33476
rect 25087 33473 25099 33507
rect 30009 33507 30067 33513
rect 30009 33504 30021 33507
rect 25041 33467 25099 33473
rect 28644 33476 30021 33504
rect 6733 33303 6791 33309
rect 6733 33269 6745 33303
rect 6779 33300 6791 33303
rect 6822 33300 6828 33312
rect 6779 33272 6828 33300
rect 6779 33269 6791 33272
rect 6733 33263 6791 33269
rect 6822 33260 6828 33272
rect 6880 33260 6886 33312
rect 7285 33303 7343 33309
rect 7285 33269 7297 33303
rect 7331 33300 7343 33303
rect 8018 33300 8024 33312
rect 7331 33272 8024 33300
rect 7331 33269 7343 33272
rect 7285 33263 7343 33269
rect 8018 33260 8024 33272
rect 8076 33260 8082 33312
rect 24394 33300 24400 33312
rect 24355 33272 24400 33300
rect 24394 33260 24400 33272
rect 24452 33260 24458 33312
rect 27338 33260 27344 33312
rect 27396 33300 27402 33312
rect 28644 33309 28672 33476
rect 30009 33473 30021 33476
rect 30055 33473 30067 33507
rect 33594 33504 33600 33516
rect 33555 33476 33600 33504
rect 30009 33467 30067 33473
rect 33594 33464 33600 33476
rect 33652 33464 33658 33516
rect 38930 33504 38936 33516
rect 38891 33476 38936 33504
rect 38930 33464 38936 33476
rect 38988 33464 38994 33516
rect 43441 33507 43499 33513
rect 43441 33473 43453 33507
rect 43487 33504 43499 33507
rect 43898 33504 43904 33516
rect 43487 33476 43904 33504
rect 43487 33473 43499 33476
rect 43441 33467 43499 33473
rect 43898 33464 43904 33476
rect 43956 33464 43962 33516
rect 48406 33504 48412 33516
rect 48367 33476 48412 33504
rect 48406 33464 48412 33476
rect 48464 33464 48470 33516
rect 52638 33464 52644 33516
rect 52696 33504 52702 33516
rect 52917 33507 52975 33513
rect 52917 33504 52929 33507
rect 52696 33476 52929 33504
rect 52696 33464 52702 33476
rect 52917 33473 52929 33476
rect 52963 33473 52975 33507
rect 52917 33467 52975 33473
rect 57149 33507 57207 33513
rect 57149 33473 57161 33507
rect 57195 33504 57207 33507
rect 57790 33504 57796 33516
rect 57195 33476 57796 33504
rect 57195 33473 57207 33476
rect 57149 33467 57207 33473
rect 57790 33464 57796 33476
rect 57848 33464 57854 33516
rect 57885 33507 57943 33513
rect 57885 33473 57897 33507
rect 57931 33473 57943 33507
rect 57885 33467 57943 33473
rect 56594 33396 56600 33448
rect 56652 33436 56658 33448
rect 57900 33436 57928 33467
rect 56652 33408 57928 33436
rect 56652 33396 56658 33408
rect 30193 33371 30251 33377
rect 30193 33337 30205 33371
rect 30239 33368 30251 33371
rect 36262 33368 36268 33380
rect 30239 33340 36268 33368
rect 30239 33337 30251 33340
rect 30193 33331 30251 33337
rect 36262 33328 36268 33340
rect 36320 33328 36326 33380
rect 58066 33368 58072 33380
rect 58027 33340 58072 33368
rect 58066 33328 58072 33340
rect 58124 33328 58130 33380
rect 28629 33303 28687 33309
rect 28629 33300 28641 33303
rect 27396 33272 28641 33300
rect 27396 33260 27402 33272
rect 28629 33269 28641 33272
rect 28675 33269 28687 33303
rect 28629 33263 28687 33269
rect 35894 33260 35900 33312
rect 35952 33300 35958 33312
rect 37553 33303 37611 33309
rect 37553 33300 37565 33303
rect 35952 33272 37565 33300
rect 35952 33260 35958 33272
rect 37553 33269 37565 33272
rect 37599 33300 37611 33303
rect 37734 33300 37740 33312
rect 37599 33272 37740 33300
rect 37599 33269 37611 33272
rect 37553 33263 37611 33269
rect 37734 33260 37740 33272
rect 37792 33260 37798 33312
rect 57333 33303 57391 33309
rect 57333 33269 57345 33303
rect 57379 33300 57391 33303
rect 57514 33300 57520 33312
rect 57379 33272 57520 33300
rect 57379 33269 57391 33272
rect 57333 33263 57391 33269
rect 57514 33260 57520 33272
rect 57572 33260 57578 33312
rect 1104 33210 58880 33232
rect 1104 33158 8174 33210
rect 8226 33158 8238 33210
rect 8290 33158 8302 33210
rect 8354 33158 8366 33210
rect 8418 33158 8430 33210
rect 8482 33158 22622 33210
rect 22674 33158 22686 33210
rect 22738 33158 22750 33210
rect 22802 33158 22814 33210
rect 22866 33158 22878 33210
rect 22930 33158 37070 33210
rect 37122 33158 37134 33210
rect 37186 33158 37198 33210
rect 37250 33158 37262 33210
rect 37314 33158 37326 33210
rect 37378 33158 51518 33210
rect 51570 33158 51582 33210
rect 51634 33158 51646 33210
rect 51698 33158 51710 33210
rect 51762 33158 51774 33210
rect 51826 33158 58880 33210
rect 1104 33136 58880 33158
rect 4525 33099 4583 33105
rect 4525 33065 4537 33099
rect 4571 33096 4583 33099
rect 4614 33096 4620 33108
rect 4571 33068 4620 33096
rect 4571 33065 4583 33068
rect 4525 33059 4583 33065
rect 4614 33056 4620 33068
rect 4672 33056 4678 33108
rect 19426 33096 19432 33108
rect 19387 33068 19432 33096
rect 19426 33056 19432 33068
rect 19484 33056 19490 33108
rect 32493 33099 32551 33105
rect 32493 33065 32505 33099
rect 32539 33096 32551 33099
rect 33594 33096 33600 33108
rect 32539 33068 33600 33096
rect 32539 33065 32551 33068
rect 32493 33059 32551 33065
rect 33594 33056 33600 33068
rect 33652 33056 33658 33108
rect 37921 33099 37979 33105
rect 37921 33065 37933 33099
rect 37967 33096 37979 33099
rect 38930 33096 38936 33108
rect 37967 33068 38936 33096
rect 37967 33065 37979 33068
rect 37921 33059 37979 33065
rect 38930 33056 38936 33068
rect 38988 33056 38994 33108
rect 57517 33099 57575 33105
rect 57517 33065 57529 33099
rect 57563 33096 57575 33099
rect 57790 33096 57796 33108
rect 57563 33068 57796 33096
rect 57563 33065 57575 33068
rect 57517 33059 57575 33065
rect 57790 33056 57796 33068
rect 57848 33056 57854 33108
rect 4341 32895 4399 32901
rect 4341 32861 4353 32895
rect 4387 32892 4399 32895
rect 4430 32892 4436 32904
rect 4387 32864 4436 32892
rect 4387 32861 4399 32864
rect 4341 32855 4399 32861
rect 4430 32852 4436 32864
rect 4488 32852 4494 32904
rect 5166 32892 5172 32904
rect 5127 32864 5172 32892
rect 5166 32852 5172 32864
rect 5224 32852 5230 32904
rect 5442 32892 5448 32904
rect 5403 32864 5448 32892
rect 5442 32852 5448 32864
rect 5500 32852 5506 32904
rect 6181 32895 6239 32901
rect 6181 32861 6193 32895
rect 6227 32892 6239 32895
rect 6546 32892 6552 32904
rect 6227 32864 6552 32892
rect 6227 32861 6239 32864
rect 6181 32855 6239 32861
rect 6546 32852 6552 32864
rect 6604 32852 6610 32904
rect 18690 32892 18696 32904
rect 18603 32864 18696 32892
rect 18690 32852 18696 32864
rect 18748 32892 18754 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 18748 32864 19257 32892
rect 18748 32852 18754 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 22925 32895 22983 32901
rect 22925 32861 22937 32895
rect 22971 32892 22983 32895
rect 32309 32895 32367 32901
rect 22971 32864 23520 32892
rect 22971 32861 22983 32864
rect 22925 32855 22983 32861
rect 5460 32824 5488 32852
rect 6825 32827 6883 32833
rect 6825 32824 6837 32827
rect 5460 32796 6837 32824
rect 6825 32793 6837 32796
rect 6871 32824 6883 32827
rect 6914 32824 6920 32836
rect 6871 32796 6920 32824
rect 6871 32793 6883 32796
rect 6825 32787 6883 32793
rect 6914 32784 6920 32796
rect 6972 32784 6978 32836
rect 6362 32756 6368 32768
rect 6323 32728 6368 32756
rect 6362 32716 6368 32728
rect 6420 32716 6426 32768
rect 7006 32716 7012 32768
rect 7064 32756 7070 32768
rect 7377 32759 7435 32765
rect 7377 32756 7389 32759
rect 7064 32728 7389 32756
rect 7064 32716 7070 32728
rect 7377 32725 7389 32728
rect 7423 32725 7435 32759
rect 7377 32719 7435 32725
rect 9398 32716 9404 32768
rect 9456 32756 9462 32768
rect 23492 32765 23520 32864
rect 32309 32861 32321 32895
rect 32355 32892 32367 32895
rect 32355 32864 32996 32892
rect 32355 32861 32367 32864
rect 32309 32855 32367 32861
rect 32968 32768 32996 32864
rect 35802 32852 35808 32904
rect 35860 32892 35866 32904
rect 36081 32895 36139 32901
rect 36081 32892 36093 32895
rect 35860 32864 36093 32892
rect 35860 32852 35866 32864
rect 36081 32861 36093 32864
rect 36127 32861 36139 32895
rect 36081 32855 36139 32861
rect 36357 32895 36415 32901
rect 36357 32861 36369 32895
rect 36403 32861 36415 32895
rect 36357 32855 36415 32861
rect 36372 32824 36400 32855
rect 36446 32852 36452 32904
rect 36504 32892 36510 32904
rect 37001 32895 37059 32901
rect 37001 32892 37013 32895
rect 36504 32864 37013 32892
rect 36504 32852 36510 32864
rect 37001 32861 37013 32864
rect 37047 32861 37059 32895
rect 37734 32892 37740 32904
rect 37695 32864 37740 32892
rect 37001 32855 37059 32861
rect 37734 32852 37740 32864
rect 37792 32852 37798 32904
rect 39853 32895 39911 32901
rect 39853 32861 39865 32895
rect 39899 32861 39911 32895
rect 39853 32855 39911 32861
rect 35866 32796 36400 32824
rect 37277 32827 37335 32833
rect 22741 32759 22799 32765
rect 22741 32756 22753 32759
rect 9456 32728 22753 32756
rect 9456 32716 9462 32728
rect 22741 32725 22753 32728
rect 22787 32725 22799 32759
rect 22741 32719 22799 32725
rect 23477 32759 23535 32765
rect 23477 32725 23489 32759
rect 23523 32756 23535 32759
rect 24302 32756 24308 32768
rect 23523 32728 24308 32756
rect 23523 32725 23535 32728
rect 23477 32719 23535 32725
rect 24302 32716 24308 32728
rect 24360 32716 24366 32768
rect 32950 32756 32956 32768
rect 32911 32728 32956 32756
rect 32950 32716 32956 32728
rect 33008 32716 33014 32768
rect 35621 32759 35679 32765
rect 35621 32725 35633 32759
rect 35667 32756 35679 32759
rect 35710 32756 35716 32768
rect 35667 32728 35716 32756
rect 35667 32725 35679 32728
rect 35621 32719 35679 32725
rect 35710 32716 35716 32728
rect 35768 32756 35774 32768
rect 35866 32756 35894 32796
rect 37277 32793 37289 32827
rect 37323 32824 37335 32827
rect 37550 32824 37556 32836
rect 37323 32796 37556 32824
rect 37323 32793 37335 32796
rect 37277 32787 37335 32793
rect 37550 32784 37556 32796
rect 37608 32824 37614 32836
rect 39868 32824 39896 32855
rect 37608 32796 39896 32824
rect 37608 32784 37614 32796
rect 35768 32728 35894 32756
rect 40037 32759 40095 32765
rect 35768 32716 35774 32728
rect 40037 32725 40049 32759
rect 40083 32756 40095 32759
rect 48406 32756 48412 32768
rect 40083 32728 48412 32756
rect 40083 32725 40095 32728
rect 40037 32719 40095 32725
rect 48406 32716 48412 32728
rect 48464 32716 48470 32768
rect 52638 32716 52644 32768
rect 52696 32756 52702 32768
rect 52733 32759 52791 32765
rect 52733 32756 52745 32759
rect 52696 32728 52745 32756
rect 52696 32716 52702 32728
rect 52733 32725 52745 32728
rect 52779 32725 52791 32759
rect 52733 32719 52791 32725
rect 1104 32666 58880 32688
rect 1104 32614 15398 32666
rect 15450 32614 15462 32666
rect 15514 32614 15526 32666
rect 15578 32614 15590 32666
rect 15642 32614 15654 32666
rect 15706 32614 29846 32666
rect 29898 32614 29910 32666
rect 29962 32614 29974 32666
rect 30026 32614 30038 32666
rect 30090 32614 30102 32666
rect 30154 32614 44294 32666
rect 44346 32614 44358 32666
rect 44410 32614 44422 32666
rect 44474 32614 44486 32666
rect 44538 32614 44550 32666
rect 44602 32614 58880 32666
rect 1104 32592 58880 32614
rect 6546 32552 6552 32564
rect 6507 32524 6552 32552
rect 6546 32512 6552 32524
rect 6604 32512 6610 32564
rect 37734 32512 37740 32564
rect 37792 32552 37798 32564
rect 38562 32552 38568 32564
rect 37792 32524 38568 32552
rect 37792 32512 37798 32524
rect 38562 32512 38568 32524
rect 38620 32552 38626 32564
rect 39117 32555 39175 32561
rect 39117 32552 39129 32555
rect 38620 32524 39129 32552
rect 38620 32512 38626 32524
rect 39117 32521 39129 32524
rect 39163 32521 39175 32555
rect 39117 32515 39175 32521
rect 3421 32487 3479 32493
rect 3421 32484 3433 32487
rect 2056 32456 3433 32484
rect 2056 32425 2084 32456
rect 3421 32453 3433 32456
rect 3467 32484 3479 32487
rect 5442 32484 5448 32496
rect 3467 32456 5448 32484
rect 3467 32453 3479 32456
rect 3421 32447 3479 32453
rect 5442 32444 5448 32456
rect 5500 32484 5506 32496
rect 5721 32487 5779 32493
rect 5721 32484 5733 32487
rect 5500 32456 5733 32484
rect 5500 32444 5506 32456
rect 5721 32453 5733 32456
rect 5767 32453 5779 32487
rect 7006 32484 7012 32496
rect 5721 32447 5779 32453
rect 6886 32456 7012 32484
rect 2041 32419 2099 32425
rect 2041 32385 2053 32419
rect 2087 32385 2099 32419
rect 2774 32416 2780 32428
rect 2735 32388 2780 32416
rect 2041 32379 2099 32385
rect 2774 32376 2780 32388
rect 2832 32376 2838 32428
rect 6365 32419 6423 32425
rect 6365 32385 6377 32419
rect 6411 32416 6423 32419
rect 6886 32416 6914 32456
rect 7006 32444 7012 32456
rect 7064 32444 7070 32496
rect 7926 32444 7932 32496
rect 7984 32444 7990 32496
rect 36262 32444 36268 32496
rect 36320 32484 36326 32496
rect 36320 32456 37964 32484
rect 36320 32444 36326 32456
rect 37936 32425 37964 32456
rect 6411 32388 6914 32416
rect 37277 32419 37335 32425
rect 6411 32385 6423 32388
rect 6365 32379 6423 32385
rect 37277 32385 37289 32419
rect 37323 32385 37335 32419
rect 37277 32379 37335 32385
rect 37921 32419 37979 32425
rect 37921 32385 37933 32419
rect 37967 32385 37979 32419
rect 37921 32379 37979 32385
rect 1762 32348 1768 32360
rect 1723 32320 1768 32348
rect 1762 32308 1768 32320
rect 1820 32308 1826 32360
rect 6914 32308 6920 32360
rect 6972 32348 6978 32360
rect 7009 32351 7067 32357
rect 7009 32348 7021 32351
rect 6972 32320 7021 32348
rect 6972 32308 6978 32320
rect 7009 32317 7021 32320
rect 7055 32317 7067 32351
rect 7009 32311 7067 32317
rect 7285 32351 7343 32357
rect 7285 32317 7297 32351
rect 7331 32348 7343 32351
rect 9030 32348 9036 32360
rect 7331 32320 8340 32348
rect 8991 32320 9036 32348
rect 7331 32317 7343 32320
rect 7285 32311 7343 32317
rect 2961 32215 3019 32221
rect 2961 32181 2973 32215
rect 3007 32212 3019 32215
rect 3050 32212 3056 32224
rect 3007 32184 3056 32212
rect 3007 32181 3019 32184
rect 2961 32175 3019 32181
rect 3050 32172 3056 32184
rect 3108 32172 3114 32224
rect 4430 32172 4436 32224
rect 4488 32212 4494 32224
rect 4617 32215 4675 32221
rect 4617 32212 4629 32215
rect 4488 32184 4629 32212
rect 4488 32172 4494 32184
rect 4617 32181 4629 32184
rect 4663 32181 4675 32215
rect 8312 32212 8340 32320
rect 9030 32308 9036 32320
rect 9088 32308 9094 32360
rect 37292 32348 37320 32379
rect 37292 32320 37964 32348
rect 37936 32224 37964 32320
rect 9585 32215 9643 32221
rect 9585 32212 9597 32215
rect 8312 32184 9597 32212
rect 4617 32175 4675 32181
rect 9585 32181 9597 32184
rect 9631 32212 9643 32215
rect 24394 32212 24400 32224
rect 9631 32184 24400 32212
rect 9631 32181 9643 32184
rect 9585 32175 9643 32181
rect 24394 32172 24400 32184
rect 24452 32172 24458 32224
rect 35710 32212 35716 32224
rect 35671 32184 35716 32212
rect 35710 32172 35716 32184
rect 35768 32172 35774 32224
rect 35802 32172 35808 32224
rect 35860 32212 35866 32224
rect 36265 32215 36323 32221
rect 36265 32212 36277 32215
rect 35860 32184 36277 32212
rect 35860 32172 35866 32184
rect 36265 32181 36277 32184
rect 36311 32181 36323 32215
rect 37458 32212 37464 32224
rect 37419 32184 37464 32212
rect 36265 32175 36323 32181
rect 37458 32172 37464 32184
rect 37516 32172 37522 32224
rect 37918 32172 37924 32224
rect 37976 32212 37982 32224
rect 38105 32215 38163 32221
rect 38105 32212 38117 32215
rect 37976 32184 38117 32212
rect 37976 32172 37982 32184
rect 38105 32181 38117 32184
rect 38151 32181 38163 32215
rect 38105 32175 38163 32181
rect 38470 32172 38476 32224
rect 38528 32212 38534 32224
rect 38565 32215 38623 32221
rect 38565 32212 38577 32215
rect 38528 32184 38577 32212
rect 38528 32172 38534 32184
rect 38565 32181 38577 32184
rect 38611 32181 38623 32215
rect 38565 32175 38623 32181
rect 1104 32122 58880 32144
rect 1104 32070 8174 32122
rect 8226 32070 8238 32122
rect 8290 32070 8302 32122
rect 8354 32070 8366 32122
rect 8418 32070 8430 32122
rect 8482 32070 22622 32122
rect 22674 32070 22686 32122
rect 22738 32070 22750 32122
rect 22802 32070 22814 32122
rect 22866 32070 22878 32122
rect 22930 32070 37070 32122
rect 37122 32070 37134 32122
rect 37186 32070 37198 32122
rect 37250 32070 37262 32122
rect 37314 32070 37326 32122
rect 37378 32070 51518 32122
rect 51570 32070 51582 32122
rect 51634 32070 51646 32122
rect 51698 32070 51710 32122
rect 51762 32070 51774 32122
rect 51826 32070 58880 32122
rect 1104 32048 58880 32070
rect 37277 32011 37335 32017
rect 37277 31977 37289 32011
rect 37323 32008 37335 32011
rect 37550 32008 37556 32020
rect 37323 31980 37556 32008
rect 37323 31977 37335 31980
rect 37277 31971 37335 31977
rect 37550 31968 37556 31980
rect 37608 32008 37614 32020
rect 37737 32011 37795 32017
rect 37737 32008 37749 32011
rect 37608 31980 37749 32008
rect 37608 31968 37614 31980
rect 37737 31977 37749 31980
rect 37783 31977 37795 32011
rect 37737 31971 37795 31977
rect 38562 31968 38568 32020
rect 38620 32008 38626 32020
rect 38620 31980 38976 32008
rect 38620 31968 38626 31980
rect 8018 31832 8024 31884
rect 8076 31872 8082 31884
rect 38948 31881 38976 31980
rect 9493 31875 9551 31881
rect 9493 31872 9505 31875
rect 8076 31844 9505 31872
rect 8076 31832 8082 31844
rect 9493 31841 9505 31844
rect 9539 31841 9551 31875
rect 9493 31835 9551 31841
rect 38933 31875 38991 31881
rect 38933 31841 38945 31875
rect 38979 31841 38991 31875
rect 38933 31835 38991 31841
rect 1762 31764 1768 31816
rect 1820 31804 1826 31816
rect 3145 31807 3203 31813
rect 3145 31804 3157 31807
rect 1820 31776 3157 31804
rect 1820 31764 1826 31776
rect 3145 31773 3157 31776
rect 3191 31804 3203 31807
rect 5166 31804 5172 31816
rect 3191 31776 5172 31804
rect 3191 31773 3203 31776
rect 3145 31767 3203 31773
rect 4632 31680 4660 31776
rect 5166 31764 5172 31776
rect 5224 31764 5230 31816
rect 5442 31804 5448 31816
rect 5403 31776 5448 31804
rect 5442 31764 5448 31776
rect 5500 31764 5506 31816
rect 6178 31804 6184 31816
rect 6139 31776 6184 31804
rect 6178 31764 6184 31776
rect 6236 31764 6242 31816
rect 6546 31764 6552 31816
rect 6604 31804 6610 31816
rect 7009 31807 7067 31813
rect 7009 31804 7021 31807
rect 6604 31776 7021 31804
rect 6604 31764 6610 31776
rect 7009 31773 7021 31776
rect 7055 31773 7067 31807
rect 7009 31767 7067 31773
rect 7745 31807 7803 31813
rect 7745 31773 7757 31807
rect 7791 31773 7803 31807
rect 35802 31804 35808 31816
rect 7745 31767 7803 31773
rect 35360 31776 35808 31804
rect 4614 31668 4620 31680
rect 4575 31640 4620 31668
rect 4614 31628 4620 31640
rect 4672 31628 4678 31680
rect 6362 31668 6368 31680
rect 6323 31640 6368 31668
rect 6362 31628 6368 31640
rect 6420 31668 6426 31680
rect 6825 31671 6883 31677
rect 6825 31668 6837 31671
rect 6420 31640 6837 31668
rect 6420 31628 6426 31640
rect 6825 31637 6837 31640
rect 6871 31637 6883 31671
rect 6825 31631 6883 31637
rect 7650 31628 7656 31680
rect 7708 31668 7714 31680
rect 7760 31668 7788 31767
rect 8941 31671 8999 31677
rect 8941 31668 8953 31671
rect 7708 31640 8953 31668
rect 7708 31628 7714 31640
rect 8941 31637 8953 31640
rect 8987 31637 8999 31671
rect 8941 31631 8999 31637
rect 35158 31628 35164 31680
rect 35216 31668 35222 31680
rect 35360 31677 35388 31776
rect 35802 31764 35808 31776
rect 35860 31804 35866 31816
rect 36081 31807 36139 31813
rect 36081 31804 36093 31807
rect 35860 31776 36093 31804
rect 35860 31764 35866 31776
rect 36081 31773 36093 31776
rect 36127 31773 36139 31807
rect 36081 31767 36139 31773
rect 36357 31807 36415 31813
rect 36357 31773 36369 31807
rect 36403 31804 36415 31807
rect 37093 31807 37151 31813
rect 36403 31776 36437 31804
rect 36403 31773 36415 31776
rect 36357 31767 36415 31773
rect 37093 31773 37105 31807
rect 37139 31804 37151 31807
rect 37458 31804 37464 31816
rect 37139 31776 37464 31804
rect 37139 31773 37151 31776
rect 37093 31767 37151 31773
rect 35710 31696 35716 31748
rect 35768 31736 35774 31748
rect 36372 31736 36400 31767
rect 37458 31764 37464 31776
rect 37516 31764 37522 31816
rect 37918 31804 37924 31816
rect 37879 31776 37924 31804
rect 37918 31764 37924 31776
rect 37976 31764 37982 31816
rect 38470 31764 38476 31816
rect 38528 31804 38534 31816
rect 38657 31807 38715 31813
rect 38657 31804 38669 31807
rect 38528 31776 38669 31804
rect 38528 31764 38534 31776
rect 38657 31773 38669 31776
rect 38703 31773 38715 31807
rect 38657 31767 38715 31773
rect 38488 31736 38516 31764
rect 35768 31708 38516 31736
rect 35768 31696 35774 31708
rect 35345 31671 35403 31677
rect 35345 31668 35357 31671
rect 35216 31640 35357 31668
rect 35216 31628 35222 31640
rect 35345 31637 35357 31640
rect 35391 31637 35403 31671
rect 35345 31631 35403 31637
rect 1104 31578 58880 31600
rect 1104 31526 15398 31578
rect 15450 31526 15462 31578
rect 15514 31526 15526 31578
rect 15578 31526 15590 31578
rect 15642 31526 15654 31578
rect 15706 31526 29846 31578
rect 29898 31526 29910 31578
rect 29962 31526 29974 31578
rect 30026 31526 30038 31578
rect 30090 31526 30102 31578
rect 30154 31526 44294 31578
rect 44346 31526 44358 31578
rect 44410 31526 44422 31578
rect 44474 31526 44486 31578
rect 44538 31526 44550 31578
rect 44602 31526 58880 31578
rect 1104 31504 58880 31526
rect 36725 31467 36783 31473
rect 36725 31433 36737 31467
rect 36771 31464 36783 31467
rect 37277 31467 37335 31473
rect 37277 31464 37289 31467
rect 36771 31436 37289 31464
rect 36771 31433 36783 31436
rect 36725 31427 36783 31433
rect 37277 31433 37289 31436
rect 37323 31464 37335 31467
rect 37550 31464 37556 31476
rect 37323 31436 37556 31464
rect 37323 31433 37335 31436
rect 37277 31427 37335 31433
rect 37550 31424 37556 31436
rect 37608 31424 37614 31476
rect 38470 31424 38476 31476
rect 38528 31464 38534 31476
rect 38933 31467 38991 31473
rect 38933 31464 38945 31467
rect 38528 31436 38945 31464
rect 38528 31424 38534 31436
rect 38933 31433 38945 31436
rect 38979 31433 38991 31467
rect 38933 31427 38991 31433
rect 3050 31356 3056 31408
rect 3108 31396 3114 31408
rect 5810 31396 5816 31408
rect 3108 31368 5816 31396
rect 3108 31356 3114 31368
rect 5810 31356 5816 31368
rect 5868 31396 5874 31408
rect 6362 31396 6368 31408
rect 5868 31368 6368 31396
rect 5868 31356 5874 31368
rect 6362 31356 6368 31368
rect 6420 31356 6426 31408
rect 38488 31396 38516 31424
rect 38212 31368 38516 31396
rect 4893 31331 4951 31337
rect 4893 31297 4905 31331
rect 4939 31328 4951 31331
rect 5442 31328 5448 31340
rect 4939 31300 5448 31328
rect 4939 31297 4951 31300
rect 4893 31291 4951 31297
rect 5442 31288 5448 31300
rect 5500 31288 5506 31340
rect 5629 31331 5687 31337
rect 5629 31297 5641 31331
rect 5675 31328 5687 31331
rect 6178 31328 6184 31340
rect 5675 31300 6184 31328
rect 5675 31297 5687 31300
rect 5629 31291 5687 31297
rect 6178 31288 6184 31300
rect 6236 31328 6242 31340
rect 6549 31331 6607 31337
rect 6549 31328 6561 31331
rect 6236 31300 6561 31328
rect 6236 31288 6242 31300
rect 6549 31297 6561 31300
rect 6595 31297 6607 31331
rect 6549 31291 6607 31297
rect 7285 31331 7343 31337
rect 7285 31297 7297 31331
rect 7331 31328 7343 31331
rect 7650 31328 7656 31340
rect 7331 31300 7656 31328
rect 7331 31297 7343 31300
rect 7285 31291 7343 31297
rect 7650 31288 7656 31300
rect 7708 31288 7714 31340
rect 35069 31331 35127 31337
rect 35069 31297 35081 31331
rect 35115 31328 35127 31331
rect 35710 31328 35716 31340
rect 35115 31300 35716 31328
rect 35115 31297 35127 31300
rect 35069 31291 35127 31297
rect 35710 31288 35716 31300
rect 35768 31328 35774 31340
rect 35805 31331 35863 31337
rect 35805 31328 35817 31331
rect 35768 31300 35817 31328
rect 35768 31288 35774 31300
rect 35805 31297 35817 31300
rect 35851 31297 35863 31331
rect 35805 31291 35863 31297
rect 36541 31331 36599 31337
rect 36541 31297 36553 31331
rect 36587 31328 36599 31331
rect 37458 31328 37464 31340
rect 36587 31300 37464 31328
rect 36587 31297 36599 31300
rect 36541 31291 36599 31297
rect 37458 31288 37464 31300
rect 37516 31288 37522 31340
rect 38212 31337 38240 31368
rect 38197 31331 38255 31337
rect 38197 31297 38209 31331
rect 38243 31297 38255 31331
rect 38197 31291 38255 31297
rect 38473 31331 38531 31337
rect 38473 31297 38485 31331
rect 38519 31328 38531 31331
rect 38562 31328 38568 31340
rect 38519 31300 38568 31328
rect 38519 31297 38531 31300
rect 38473 31291 38531 31297
rect 38562 31288 38568 31300
rect 38620 31328 38626 31340
rect 39485 31331 39543 31337
rect 39485 31328 39497 31331
rect 38620 31300 39497 31328
rect 38620 31288 38626 31300
rect 39485 31297 39497 31300
rect 39531 31297 39543 31331
rect 45830 31328 45836 31340
rect 45791 31300 45836 31328
rect 39485 31291 39543 31297
rect 45830 31288 45836 31300
rect 45888 31328 45894 31340
rect 46477 31331 46535 31337
rect 46477 31328 46489 31331
rect 45888 31300 46489 31328
rect 45888 31288 45894 31300
rect 46477 31297 46489 31300
rect 46523 31297 46535 31331
rect 46477 31291 46535 31297
rect 4617 31263 4675 31269
rect 4617 31229 4629 31263
rect 4663 31229 4675 31263
rect 4617 31223 4675 31229
rect 7561 31263 7619 31269
rect 7561 31229 7573 31263
rect 7607 31260 7619 31263
rect 8018 31260 8024 31272
rect 7607 31232 8024 31260
rect 7607 31229 7619 31232
rect 7561 31223 7619 31229
rect 4632 31136 4660 31223
rect 8018 31220 8024 31232
rect 8076 31260 8082 31272
rect 8573 31263 8631 31269
rect 8573 31260 8585 31263
rect 8076 31232 8585 31260
rect 8076 31220 8082 31232
rect 8573 31229 8585 31232
rect 8619 31229 8631 31263
rect 8573 31223 8631 31229
rect 35158 31220 35164 31272
rect 35216 31260 35222 31272
rect 35529 31263 35587 31269
rect 35529 31260 35541 31263
rect 35216 31232 35541 31260
rect 35216 31220 35222 31232
rect 35529 31229 35541 31232
rect 35575 31229 35587 31263
rect 35529 31223 35587 31229
rect 46017 31195 46075 31201
rect 46017 31161 46029 31195
rect 46063 31192 46075 31195
rect 46063 31164 55214 31192
rect 46063 31161 46075 31164
rect 46017 31155 46075 31161
rect 4157 31127 4215 31133
rect 4157 31093 4169 31127
rect 4203 31124 4215 31127
rect 4614 31124 4620 31136
rect 4203 31096 4620 31124
rect 4203 31093 4215 31096
rect 4157 31087 4215 31093
rect 4614 31084 4620 31096
rect 4672 31084 4678 31136
rect 7650 31084 7656 31136
rect 7708 31124 7714 31136
rect 8021 31127 8079 31133
rect 8021 31124 8033 31127
rect 7708 31096 8033 31124
rect 7708 31084 7714 31096
rect 8021 31093 8033 31096
rect 8067 31093 8079 31127
rect 55186 31124 55214 31164
rect 56594 31124 56600 31136
rect 55186 31096 56600 31124
rect 8021 31087 8079 31093
rect 56594 31084 56600 31096
rect 56652 31084 56658 31136
rect 1104 31034 58880 31056
rect 1104 30982 8174 31034
rect 8226 30982 8238 31034
rect 8290 30982 8302 31034
rect 8354 30982 8366 31034
rect 8418 30982 8430 31034
rect 8482 30982 22622 31034
rect 22674 30982 22686 31034
rect 22738 30982 22750 31034
rect 22802 30982 22814 31034
rect 22866 30982 22878 31034
rect 22930 30982 37070 31034
rect 37122 30982 37134 31034
rect 37186 30982 37198 31034
rect 37250 30982 37262 31034
rect 37314 30982 37326 31034
rect 37378 30982 51518 31034
rect 51570 30982 51582 31034
rect 51634 30982 51646 31034
rect 51698 30982 51710 31034
rect 51762 30982 51774 31034
rect 51826 30982 58880 31034
rect 1104 30960 58880 30982
rect 1670 30880 1676 30932
rect 1728 30920 1734 30932
rect 2225 30923 2283 30929
rect 2225 30920 2237 30923
rect 1728 30892 2237 30920
rect 1728 30880 1734 30892
rect 2225 30889 2237 30892
rect 2271 30889 2283 30923
rect 2225 30883 2283 30889
rect 5810 30880 5816 30932
rect 5868 30920 5874 30932
rect 6365 30923 6423 30929
rect 6365 30920 6377 30923
rect 5868 30892 6377 30920
rect 5868 30880 5874 30892
rect 6365 30889 6377 30892
rect 6411 30920 6423 30923
rect 6822 30920 6828 30932
rect 6411 30892 6828 30920
rect 6411 30889 6423 30892
rect 6365 30883 6423 30889
rect 6822 30880 6828 30892
rect 6880 30880 6886 30932
rect 37277 30923 37335 30929
rect 37277 30889 37289 30923
rect 37323 30920 37335 30923
rect 37550 30920 37556 30932
rect 37323 30892 37556 30920
rect 37323 30889 37335 30892
rect 37277 30883 37335 30889
rect 37550 30880 37556 30892
rect 37608 30920 37614 30932
rect 37737 30923 37795 30929
rect 37737 30920 37749 30923
rect 37608 30892 37749 30920
rect 37608 30880 37614 30892
rect 37737 30889 37749 30892
rect 37783 30889 37795 30923
rect 37737 30883 37795 30889
rect 38562 30880 38568 30932
rect 38620 30920 38626 30932
rect 38620 30892 38884 30920
rect 38620 30880 38626 30892
rect 38856 30852 38884 30892
rect 38856 30824 38976 30852
rect 38948 30793 38976 30824
rect 38933 30787 38991 30793
rect 38933 30753 38945 30787
rect 38979 30753 38991 30787
rect 38933 30747 38991 30753
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30685 1731 30719
rect 1673 30679 1731 30685
rect 2409 30719 2467 30725
rect 2409 30685 2421 30719
rect 2455 30716 2467 30719
rect 2866 30716 2872 30728
rect 2455 30688 2872 30716
rect 2455 30685 2467 30688
rect 2409 30679 2467 30685
rect 1688 30648 1716 30679
rect 2866 30676 2872 30688
rect 2924 30676 2930 30728
rect 3050 30716 3056 30728
rect 3011 30688 3056 30716
rect 3050 30676 3056 30688
rect 3108 30676 3114 30728
rect 4614 30676 4620 30728
rect 4672 30716 4678 30728
rect 5169 30719 5227 30725
rect 5169 30716 5181 30719
rect 4672 30688 5181 30716
rect 4672 30676 4678 30688
rect 5169 30685 5181 30688
rect 5215 30685 5227 30719
rect 5442 30716 5448 30728
rect 5403 30688 5448 30716
rect 5169 30679 5227 30685
rect 5442 30676 5448 30688
rect 5500 30676 5506 30728
rect 6178 30716 6184 30728
rect 6139 30688 6184 30716
rect 6178 30676 6184 30688
rect 6236 30676 6242 30728
rect 6546 30676 6552 30728
rect 6604 30716 6610 30728
rect 7009 30719 7067 30725
rect 7009 30716 7021 30719
rect 6604 30688 7021 30716
rect 6604 30676 6610 30688
rect 7009 30685 7021 30688
rect 7055 30685 7067 30719
rect 7009 30679 7067 30685
rect 7745 30719 7803 30725
rect 7745 30685 7757 30719
rect 7791 30685 7803 30719
rect 8018 30716 8024 30728
rect 7979 30688 8024 30716
rect 7745 30679 7803 30685
rect 1688 30620 2912 30648
rect 1486 30580 1492 30592
rect 1447 30552 1492 30580
rect 1486 30540 1492 30552
rect 1544 30540 1550 30592
rect 2884 30589 2912 30620
rect 2869 30583 2927 30589
rect 2869 30549 2881 30583
rect 2915 30549 2927 30583
rect 4614 30580 4620 30592
rect 4575 30552 4620 30580
rect 2869 30543 2927 30549
rect 4614 30540 4620 30552
rect 4672 30540 4678 30592
rect 7650 30540 7656 30592
rect 7708 30580 7714 30592
rect 7760 30580 7788 30679
rect 8018 30676 8024 30688
rect 8076 30676 8082 30728
rect 35802 30676 35808 30728
rect 35860 30716 35866 30728
rect 36081 30719 36139 30725
rect 36081 30716 36093 30719
rect 35860 30688 36093 30716
rect 35860 30676 35866 30688
rect 36081 30685 36093 30688
rect 36127 30685 36139 30719
rect 36081 30679 36139 30685
rect 36357 30719 36415 30725
rect 36357 30685 36369 30719
rect 36403 30685 36415 30719
rect 36357 30679 36415 30685
rect 37093 30719 37151 30725
rect 37093 30685 37105 30719
rect 37139 30716 37151 30719
rect 37458 30716 37464 30728
rect 37139 30688 37464 30716
rect 37139 30685 37151 30688
rect 37093 30679 37151 30685
rect 36372 30648 36400 30679
rect 37458 30676 37464 30688
rect 37516 30676 37522 30728
rect 37918 30716 37924 30728
rect 37879 30688 37924 30716
rect 37918 30676 37924 30688
rect 37976 30676 37982 30728
rect 38470 30676 38476 30728
rect 38528 30716 38534 30728
rect 38657 30719 38715 30725
rect 38657 30716 38669 30719
rect 38528 30688 38669 30716
rect 38528 30676 38534 30688
rect 38657 30685 38669 30688
rect 38703 30685 38715 30719
rect 38657 30679 38715 30685
rect 37366 30648 37372 30660
rect 35866 30620 37372 30648
rect 8941 30583 8999 30589
rect 8941 30580 8953 30583
rect 7708 30552 8953 30580
rect 7708 30540 7714 30552
rect 8941 30549 8953 30552
rect 8987 30549 8999 30583
rect 8941 30543 8999 30549
rect 35069 30583 35127 30589
rect 35069 30549 35081 30583
rect 35115 30580 35127 30583
rect 35158 30580 35164 30592
rect 35115 30552 35164 30580
rect 35115 30549 35127 30552
rect 35069 30543 35127 30549
rect 35158 30540 35164 30552
rect 35216 30540 35222 30592
rect 35342 30540 35348 30592
rect 35400 30580 35406 30592
rect 35529 30583 35587 30589
rect 35529 30580 35541 30583
rect 35400 30552 35541 30580
rect 35400 30540 35406 30552
rect 35529 30549 35541 30552
rect 35575 30580 35587 30583
rect 35866 30580 35894 30620
rect 37366 30608 37372 30620
rect 37424 30608 37430 30660
rect 35575 30552 35894 30580
rect 35575 30549 35587 30552
rect 35529 30543 35587 30549
rect 1104 30490 58880 30512
rect 1104 30438 15398 30490
rect 15450 30438 15462 30490
rect 15514 30438 15526 30490
rect 15578 30438 15590 30490
rect 15642 30438 15654 30490
rect 15706 30438 29846 30490
rect 29898 30438 29910 30490
rect 29962 30438 29974 30490
rect 30026 30438 30038 30490
rect 30090 30438 30102 30490
rect 30154 30438 44294 30490
rect 44346 30438 44358 30490
rect 44410 30438 44422 30490
rect 44474 30438 44486 30490
rect 44538 30438 44550 30490
rect 44602 30438 58880 30490
rect 1104 30416 58880 30438
rect 5810 30376 5816 30388
rect 5771 30348 5816 30376
rect 5810 30336 5816 30348
rect 5868 30336 5874 30388
rect 6178 30336 6184 30388
rect 6236 30376 6242 30388
rect 6549 30379 6607 30385
rect 6549 30376 6561 30379
rect 6236 30348 6561 30376
rect 6236 30336 6242 30348
rect 6549 30345 6561 30348
rect 6595 30345 6607 30379
rect 6549 30339 6607 30345
rect 37366 30336 37372 30388
rect 37424 30376 37430 30388
rect 37461 30379 37519 30385
rect 37461 30376 37473 30379
rect 37424 30348 37473 30376
rect 37424 30336 37430 30348
rect 37461 30345 37473 30348
rect 37507 30376 37519 30379
rect 38470 30376 38476 30388
rect 37507 30348 38476 30376
rect 37507 30345 37519 30348
rect 37461 30339 37519 30345
rect 38470 30336 38476 30348
rect 38528 30336 38534 30388
rect 7006 30308 7012 30320
rect 5644 30280 7012 30308
rect 4893 30243 4951 30249
rect 4893 30209 4905 30243
rect 4939 30240 4951 30243
rect 5442 30240 5448 30252
rect 4939 30212 5448 30240
rect 4939 30209 4951 30212
rect 4893 30203 4951 30209
rect 5442 30200 5448 30212
rect 5500 30200 5506 30252
rect 5644 30249 5672 30280
rect 7006 30268 7012 30280
rect 7064 30268 7070 30320
rect 5629 30243 5687 30249
rect 5629 30209 5641 30243
rect 5675 30209 5687 30243
rect 5629 30203 5687 30209
rect 6365 30243 6423 30249
rect 6365 30209 6377 30243
rect 6411 30240 6423 30243
rect 6546 30240 6552 30252
rect 6411 30212 6552 30240
rect 6411 30209 6423 30212
rect 6365 30203 6423 30209
rect 6546 30200 6552 30212
rect 6604 30200 6610 30252
rect 6822 30200 6828 30252
rect 6880 30240 6886 30252
rect 7834 30240 7840 30252
rect 6880 30212 7840 30240
rect 6880 30200 6886 30212
rect 7834 30200 7840 30212
rect 7892 30200 7898 30252
rect 14366 30200 14372 30252
rect 14424 30240 14430 30252
rect 14921 30243 14979 30249
rect 14921 30240 14933 30243
rect 14424 30212 14933 30240
rect 14424 30200 14430 30212
rect 14921 30209 14933 30212
rect 14967 30209 14979 30243
rect 19518 30240 19524 30252
rect 19479 30212 19524 30240
rect 14921 30203 14979 30209
rect 19518 30200 19524 30212
rect 19576 30200 19582 30252
rect 4614 30172 4620 30184
rect 4172 30144 4620 30172
rect 4172 30048 4200 30144
rect 4614 30132 4620 30144
rect 4672 30132 4678 30184
rect 5460 30104 5488 30200
rect 14550 30132 14556 30184
rect 14608 30172 14614 30184
rect 14829 30175 14887 30181
rect 14829 30172 14841 30175
rect 14608 30144 14841 30172
rect 14608 30132 14614 30144
rect 14829 30141 14841 30144
rect 14875 30141 14887 30175
rect 14829 30135 14887 30141
rect 35989 30107 36047 30113
rect 5460 30076 7144 30104
rect 4154 30036 4160 30048
rect 4115 30008 4160 30036
rect 4154 29996 4160 30008
rect 4212 29996 4218 30048
rect 7116 30045 7144 30076
rect 35989 30073 36001 30107
rect 36035 30104 36047 30107
rect 37921 30107 37979 30113
rect 37921 30104 37933 30107
rect 36035 30076 37933 30104
rect 36035 30073 36047 30076
rect 35989 30067 36047 30073
rect 37921 30073 37933 30076
rect 37967 30073 37979 30107
rect 37921 30067 37979 30073
rect 7101 30039 7159 30045
rect 7101 30005 7113 30039
rect 7147 30036 7159 30039
rect 7650 30036 7656 30048
rect 7147 30008 7656 30036
rect 7147 30005 7159 30008
rect 7101 29999 7159 30005
rect 7650 29996 7656 30008
rect 7708 29996 7714 30048
rect 8018 29996 8024 30048
rect 8076 30036 8082 30048
rect 8113 30039 8171 30045
rect 8113 30036 8125 30039
rect 8076 30008 8125 30036
rect 8076 29996 8082 30008
rect 8113 30005 8125 30008
rect 8159 30005 8171 30039
rect 15194 30036 15200 30048
rect 15155 30008 15200 30036
rect 8113 29999 8171 30005
rect 15194 29996 15200 30008
rect 15252 29996 15258 30048
rect 19521 30039 19579 30045
rect 19521 30005 19533 30039
rect 19567 30036 19579 30039
rect 20714 30036 20720 30048
rect 19567 30008 20720 30036
rect 19567 30005 19579 30008
rect 19521 29999 19579 30005
rect 20714 29996 20720 30008
rect 20772 29996 20778 30048
rect 35802 29996 35808 30048
rect 35860 30036 35866 30048
rect 36004 30036 36032 30067
rect 35860 30008 36032 30036
rect 35860 29996 35866 30008
rect 1104 29946 58880 29968
rect 1104 29894 8174 29946
rect 8226 29894 8238 29946
rect 8290 29894 8302 29946
rect 8354 29894 8366 29946
rect 8418 29894 8430 29946
rect 8482 29894 22622 29946
rect 22674 29894 22686 29946
rect 22738 29894 22750 29946
rect 22802 29894 22814 29946
rect 22866 29894 22878 29946
rect 22930 29894 37070 29946
rect 37122 29894 37134 29946
rect 37186 29894 37198 29946
rect 37250 29894 37262 29946
rect 37314 29894 37326 29946
rect 37378 29894 51518 29946
rect 51570 29894 51582 29946
rect 51634 29894 51646 29946
rect 51698 29894 51710 29946
rect 51762 29894 51774 29946
rect 51826 29894 58880 29946
rect 1104 29872 58880 29894
rect 15194 29792 15200 29844
rect 15252 29832 15258 29844
rect 37277 29835 37335 29841
rect 15252 29804 22094 29832
rect 15252 29792 15258 29804
rect 6914 29764 6920 29776
rect 5092 29736 6920 29764
rect 2498 29656 2504 29708
rect 2556 29696 2562 29708
rect 3237 29699 3295 29705
rect 3237 29696 3249 29699
rect 2556 29668 3249 29696
rect 2556 29656 2562 29668
rect 3237 29665 3249 29668
rect 3283 29696 3295 29699
rect 3789 29699 3847 29705
rect 3789 29696 3801 29699
rect 3283 29668 3801 29696
rect 3283 29665 3295 29668
rect 3237 29659 3295 29665
rect 3789 29665 3801 29668
rect 3835 29696 3847 29699
rect 5092 29696 5120 29736
rect 6914 29724 6920 29736
rect 6972 29724 6978 29776
rect 15013 29767 15071 29773
rect 15013 29733 15025 29767
rect 15059 29733 15071 29767
rect 15013 29727 15071 29733
rect 7009 29699 7067 29705
rect 7009 29696 7021 29699
rect 3835 29668 5120 29696
rect 5184 29668 7021 29696
rect 3835 29665 3847 29668
rect 3789 29659 3847 29665
rect 4062 29560 4068 29572
rect 4023 29532 4068 29560
rect 4062 29520 4068 29532
rect 4120 29520 4126 29572
rect 4172 29532 4554 29560
rect 3234 29452 3240 29504
rect 3292 29492 3298 29504
rect 4172 29492 4200 29532
rect 3292 29464 4200 29492
rect 4448 29492 4476 29532
rect 5184 29492 5212 29668
rect 7009 29665 7021 29668
rect 7055 29665 7067 29699
rect 14550 29696 14556 29708
rect 14511 29668 14556 29696
rect 7009 29659 7067 29665
rect 14550 29656 14556 29668
rect 14608 29656 14614 29708
rect 15028 29696 15056 29727
rect 16209 29699 16267 29705
rect 16209 29696 16221 29699
rect 15028 29668 16221 29696
rect 16209 29665 16221 29668
rect 16255 29665 16267 29699
rect 16209 29659 16267 29665
rect 17957 29699 18015 29705
rect 17957 29665 17969 29699
rect 18003 29696 18015 29699
rect 19518 29696 19524 29708
rect 18003 29668 19524 29696
rect 18003 29665 18015 29668
rect 17957 29659 18015 29665
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 20714 29696 20720 29708
rect 20675 29668 20720 29696
rect 20714 29656 20720 29668
rect 20772 29656 20778 29708
rect 22066 29696 22094 29804
rect 37277 29801 37289 29835
rect 37323 29832 37335 29835
rect 37550 29832 37556 29844
rect 37323 29804 37556 29832
rect 37323 29801 37335 29804
rect 37277 29795 37335 29801
rect 37550 29792 37556 29804
rect 37608 29792 37614 29844
rect 26881 29699 26939 29705
rect 26881 29696 26893 29699
rect 22066 29668 26893 29696
rect 26881 29665 26893 29668
rect 26927 29665 26939 29699
rect 26881 29659 26939 29665
rect 27522 29656 27528 29708
rect 27580 29696 27586 29708
rect 28629 29699 28687 29705
rect 28629 29696 28641 29699
rect 27580 29668 28641 29696
rect 27580 29656 27586 29668
rect 28629 29665 28641 29668
rect 28675 29665 28687 29699
rect 28629 29659 28687 29665
rect 5994 29628 6000 29640
rect 5955 29600 6000 29628
rect 5994 29588 6000 29600
rect 6052 29588 6058 29640
rect 14366 29588 14372 29640
rect 14424 29628 14430 29640
rect 14645 29631 14703 29637
rect 14645 29628 14657 29631
rect 14424 29600 14657 29628
rect 14424 29588 14430 29600
rect 14645 29597 14657 29600
rect 14691 29597 14703 29631
rect 14645 29591 14703 29597
rect 20993 29631 21051 29637
rect 20993 29597 21005 29631
rect 21039 29628 21051 29631
rect 24118 29628 24124 29640
rect 21039 29600 24124 29628
rect 21039 29597 21051 29600
rect 20993 29591 21051 29597
rect 7006 29520 7012 29572
rect 7064 29560 7070 29572
rect 7193 29563 7251 29569
rect 7193 29560 7205 29563
rect 7064 29532 7205 29560
rect 7064 29520 7070 29532
rect 7193 29529 7205 29532
rect 7239 29529 7251 29563
rect 16482 29560 16488 29572
rect 16443 29532 16488 29560
rect 7193 29523 7251 29529
rect 16482 29520 16488 29532
rect 16540 29520 16546 29572
rect 18598 29560 18604 29572
rect 16868 29532 16974 29560
rect 17880 29532 18604 29560
rect 4448 29464 5212 29492
rect 3292 29452 3298 29464
rect 5350 29452 5356 29504
rect 5408 29492 5414 29504
rect 5537 29495 5595 29501
rect 5537 29492 5549 29495
rect 5408 29464 5549 29492
rect 5408 29452 5414 29464
rect 5537 29461 5549 29464
rect 5583 29461 5595 29495
rect 5537 29455 5595 29461
rect 6181 29495 6239 29501
rect 6181 29461 6193 29495
rect 6227 29492 6239 29495
rect 6270 29492 6276 29504
rect 6227 29464 6276 29492
rect 6227 29461 6239 29464
rect 6181 29455 6239 29461
rect 6270 29452 6276 29464
rect 6328 29452 6334 29504
rect 8018 29452 8024 29504
rect 8076 29492 8082 29504
rect 8297 29495 8355 29501
rect 8297 29492 8309 29495
rect 8076 29464 8309 29492
rect 8076 29452 8082 29464
rect 8297 29461 8309 29464
rect 8343 29492 8355 29495
rect 9582 29492 9588 29504
rect 8343 29464 9588 29492
rect 8343 29461 8355 29464
rect 8297 29455 8355 29461
rect 9582 29452 9588 29464
rect 9640 29452 9646 29504
rect 15746 29492 15752 29504
rect 15707 29464 15752 29492
rect 15746 29452 15752 29464
rect 15804 29492 15810 29504
rect 16868 29492 16896 29532
rect 17880 29492 17908 29532
rect 18598 29520 18604 29532
rect 18656 29560 18662 29572
rect 18656 29532 19550 29560
rect 18656 29520 18662 29532
rect 20622 29520 20628 29572
rect 20680 29560 20686 29572
rect 21008 29560 21036 29591
rect 24118 29588 24124 29600
rect 24176 29588 24182 29640
rect 35158 29588 35164 29640
rect 35216 29628 35222 29640
rect 35802 29628 35808 29640
rect 35216 29600 35808 29628
rect 35216 29588 35222 29600
rect 35802 29588 35808 29600
rect 35860 29628 35866 29640
rect 36081 29631 36139 29637
rect 36081 29628 36093 29631
rect 35860 29600 36093 29628
rect 35860 29588 35866 29600
rect 36081 29597 36093 29600
rect 36127 29597 36139 29631
rect 36081 29591 36139 29597
rect 36357 29631 36415 29637
rect 36357 29597 36369 29631
rect 36403 29597 36415 29631
rect 36357 29591 36415 29597
rect 37093 29631 37151 29637
rect 37093 29597 37105 29631
rect 37139 29628 37151 29631
rect 37918 29628 37924 29640
rect 37139 29600 37924 29628
rect 37139 29597 37151 29600
rect 37093 29591 37151 29597
rect 27154 29560 27160 29572
rect 20680 29532 21036 29560
rect 27115 29532 27160 29560
rect 20680 29520 20686 29532
rect 27154 29520 27160 29532
rect 27212 29520 27218 29572
rect 36372 29560 36400 29591
rect 37918 29588 37924 29600
rect 37976 29588 37982 29640
rect 28382 29532 29684 29560
rect 19242 29492 19248 29504
rect 15804 29464 17908 29492
rect 19203 29464 19248 29492
rect 15804 29452 15810 29464
rect 19242 29452 19248 29464
rect 19300 29452 19306 29504
rect 26418 29492 26424 29504
rect 26331 29464 26424 29492
rect 26418 29452 26424 29464
rect 26476 29492 26482 29504
rect 28460 29492 28488 29532
rect 29656 29501 29684 29532
rect 35866 29532 36400 29560
rect 26476 29464 28488 29492
rect 29641 29495 29699 29501
rect 26476 29452 26482 29464
rect 29641 29461 29653 29495
rect 29687 29492 29699 29495
rect 30190 29492 30196 29504
rect 29687 29464 30196 29492
rect 29687 29461 29699 29464
rect 29641 29455 29699 29461
rect 30190 29452 30196 29464
rect 30248 29452 30254 29504
rect 35342 29452 35348 29504
rect 35400 29492 35406 29504
rect 35529 29495 35587 29501
rect 35529 29492 35541 29495
rect 35400 29464 35541 29492
rect 35400 29452 35406 29464
rect 35529 29461 35541 29464
rect 35575 29492 35587 29495
rect 35866 29492 35894 29532
rect 35575 29464 35894 29492
rect 35575 29461 35587 29464
rect 35529 29455 35587 29461
rect 1104 29402 58880 29424
rect 1104 29350 15398 29402
rect 15450 29350 15462 29402
rect 15514 29350 15526 29402
rect 15578 29350 15590 29402
rect 15642 29350 15654 29402
rect 15706 29350 29846 29402
rect 29898 29350 29910 29402
rect 29962 29350 29974 29402
rect 30026 29350 30038 29402
rect 30090 29350 30102 29402
rect 30154 29350 44294 29402
rect 44346 29350 44358 29402
rect 44410 29350 44422 29402
rect 44474 29350 44486 29402
rect 44538 29350 44550 29402
rect 44602 29350 58880 29402
rect 1104 29328 58880 29350
rect 4062 29248 4068 29300
rect 4120 29288 4126 29300
rect 4249 29291 4307 29297
rect 4249 29288 4261 29291
rect 4120 29260 4261 29288
rect 4120 29248 4126 29260
rect 4249 29257 4261 29260
rect 4295 29257 4307 29291
rect 4249 29251 4307 29257
rect 7006 29248 7012 29300
rect 7064 29248 7070 29300
rect 16482 29248 16488 29300
rect 16540 29288 16546 29300
rect 17589 29291 17647 29297
rect 17589 29288 17601 29291
rect 16540 29260 17601 29288
rect 16540 29248 16546 29260
rect 17589 29257 17601 29260
rect 17635 29257 17647 29291
rect 24118 29288 24124 29300
rect 24079 29260 24124 29288
rect 17589 29251 17647 29257
rect 24118 29248 24124 29260
rect 24176 29248 24182 29300
rect 2774 29180 2780 29232
rect 2832 29220 2838 29232
rect 3234 29220 3240 29232
rect 2832 29192 3240 29220
rect 2832 29180 2838 29192
rect 3234 29180 3240 29192
rect 3292 29180 3298 29232
rect 4154 29180 4160 29232
rect 4212 29220 4218 29232
rect 6730 29220 6736 29232
rect 4212 29192 6736 29220
rect 4212 29180 4218 29192
rect 6730 29180 6736 29192
rect 6788 29180 6794 29232
rect 7024 29220 7052 29248
rect 7024 29192 7130 29220
rect 2041 29155 2099 29161
rect 2041 29121 2053 29155
rect 2087 29152 2099 29155
rect 2498 29152 2504 29164
rect 2087 29124 2504 29152
rect 2087 29121 2099 29124
rect 2041 29115 2099 29121
rect 2498 29112 2504 29124
rect 2556 29112 2562 29164
rect 8573 29155 8631 29161
rect 8573 29121 8585 29155
rect 8619 29121 8631 29155
rect 8573 29115 8631 29121
rect 17681 29155 17739 29161
rect 17681 29121 17693 29155
rect 17727 29152 17739 29155
rect 19242 29152 19248 29164
rect 17727 29124 19248 29152
rect 17727 29121 17739 29124
rect 17681 29115 17739 29121
rect 4985 29087 5043 29093
rect 4985 29053 4997 29087
rect 5031 29053 5043 29087
rect 4985 29047 5043 29053
rect 6365 29087 6423 29093
rect 6365 29053 6377 29087
rect 6411 29084 6423 29087
rect 7006 29084 7012 29096
rect 6411 29056 7012 29084
rect 6411 29053 6423 29056
rect 6365 29047 6423 29053
rect 5000 28960 5028 29047
rect 7006 29044 7012 29056
rect 7064 29084 7070 29096
rect 8018 29084 8024 29096
rect 7064 29056 8024 29084
rect 7064 29044 7070 29056
rect 8018 29044 8024 29056
rect 8076 29044 8082 29096
rect 8113 29087 8171 29093
rect 8113 29053 8125 29087
rect 8159 29084 8171 29087
rect 8588 29084 8616 29115
rect 19242 29112 19248 29124
rect 19300 29152 19306 29164
rect 19981 29155 20039 29161
rect 19981 29152 19993 29155
rect 19300 29124 19993 29152
rect 19300 29112 19306 29124
rect 19981 29121 19993 29124
rect 20027 29121 20039 29155
rect 24136 29152 24164 29248
rect 26418 29220 26424 29232
rect 26174 29192 26424 29220
rect 26418 29180 26424 29192
rect 26476 29180 26482 29232
rect 24673 29155 24731 29161
rect 24673 29152 24685 29155
rect 24136 29124 24685 29152
rect 19981 29115 20039 29121
rect 24673 29121 24685 29124
rect 24719 29121 24731 29155
rect 26786 29152 26792 29164
rect 24673 29115 24731 29121
rect 26436 29124 26792 29152
rect 8159 29056 8616 29084
rect 8159 29053 8171 29056
rect 8113 29047 8171 29053
rect 19518 29044 19524 29096
rect 19576 29084 19582 29096
rect 19889 29087 19947 29093
rect 19889 29084 19901 29087
rect 19576 29056 19901 29084
rect 19576 29044 19582 29056
rect 19889 29053 19901 29056
rect 19935 29053 19947 29087
rect 19889 29047 19947 29053
rect 20809 29087 20867 29093
rect 20809 29053 20821 29087
rect 20855 29084 20867 29087
rect 21726 29084 21732 29096
rect 20855 29056 21732 29084
rect 20855 29053 20867 29056
rect 20809 29047 20867 29053
rect 21726 29044 21732 29056
rect 21784 29044 21790 29096
rect 26436 29093 26464 29124
rect 26786 29112 26792 29124
rect 26844 29152 26850 29164
rect 27341 29155 27399 29161
rect 27341 29152 27353 29155
rect 26844 29124 27353 29152
rect 26844 29112 26850 29124
rect 27341 29121 27353 29124
rect 27387 29121 27399 29155
rect 36262 29152 36268 29164
rect 36223 29124 36268 29152
rect 27341 29115 27399 29121
rect 36262 29112 36268 29124
rect 36320 29112 36326 29164
rect 26421 29087 26479 29093
rect 26421 29053 26433 29087
rect 26467 29053 26479 29087
rect 27522 29084 27528 29096
rect 27483 29056 27528 29084
rect 26421 29047 26479 29053
rect 27522 29044 27528 29056
rect 27580 29044 27586 29096
rect 28169 29087 28227 29093
rect 28169 29053 28181 29087
rect 28215 29084 28227 29087
rect 28902 29084 28908 29096
rect 28215 29056 28908 29084
rect 28215 29053 28227 29056
rect 28169 29047 28227 29053
rect 28902 29044 28908 29056
rect 28960 29044 28966 29096
rect 5350 29016 5356 29028
rect 5311 28988 5356 29016
rect 5350 28976 5356 28988
rect 5408 28976 5414 29028
rect 5445 29019 5503 29025
rect 5445 28985 5457 29019
rect 5491 29016 5503 29019
rect 6178 29016 6184 29028
rect 5491 28988 6184 29016
rect 5491 28985 5503 28988
rect 5445 28979 5503 28985
rect 6178 28976 6184 28988
rect 6236 28976 6242 29028
rect 8754 29016 8760 29028
rect 8715 28988 8760 29016
rect 8754 28976 8760 28988
rect 8812 28976 8818 29028
rect 36078 29016 36084 29028
rect 36039 28988 36084 29016
rect 36078 28976 36084 28988
rect 36136 28976 36142 29028
rect 2314 28908 2320 28960
rect 2372 28948 2378 28960
rect 2758 28951 2816 28957
rect 2758 28948 2770 28951
rect 2372 28920 2770 28948
rect 2372 28908 2378 28920
rect 2758 28917 2770 28920
rect 2804 28948 2816 28951
rect 4982 28948 4988 28960
rect 2804 28920 4988 28948
rect 2804 28917 2816 28920
rect 2758 28911 2816 28917
rect 4982 28908 4988 28920
rect 5040 28908 5046 28960
rect 6362 28908 6368 28960
rect 6420 28948 6426 28960
rect 6622 28951 6680 28957
rect 6622 28948 6634 28951
rect 6420 28920 6634 28948
rect 6420 28908 6426 28920
rect 6622 28917 6634 28920
rect 6668 28917 6680 28951
rect 6622 28911 6680 28917
rect 18046 28908 18052 28960
rect 18104 28948 18110 28960
rect 18877 28951 18935 28957
rect 18877 28948 18889 28951
rect 18104 28920 18889 28948
rect 18104 28908 18110 28920
rect 18877 28917 18889 28920
rect 18923 28917 18935 28951
rect 18877 28911 18935 28917
rect 24936 28951 24994 28957
rect 24936 28917 24948 28951
rect 24982 28948 24994 28951
rect 27430 28948 27436 28960
rect 24982 28920 27436 28948
rect 24982 28917 24994 28920
rect 24936 28911 24994 28917
rect 27430 28908 27436 28920
rect 27488 28908 27494 28960
rect 34790 28948 34796 28960
rect 34751 28920 34796 28948
rect 34790 28908 34796 28920
rect 34848 28908 34854 28960
rect 1104 28858 58880 28880
rect 1104 28806 8174 28858
rect 8226 28806 8238 28858
rect 8290 28806 8302 28858
rect 8354 28806 8366 28858
rect 8418 28806 8430 28858
rect 8482 28806 22622 28858
rect 22674 28806 22686 28858
rect 22738 28806 22750 28858
rect 22802 28806 22814 28858
rect 22866 28806 22878 28858
rect 22930 28806 37070 28858
rect 37122 28806 37134 28858
rect 37186 28806 37198 28858
rect 37250 28806 37262 28858
rect 37314 28806 37326 28858
rect 37378 28806 51518 28858
rect 51570 28806 51582 28858
rect 51634 28806 51646 28858
rect 51698 28806 51710 28858
rect 51762 28806 51774 28858
rect 51826 28806 58880 28858
rect 1104 28784 58880 28806
rect 5537 28747 5595 28753
rect 5537 28713 5549 28747
rect 5583 28744 5595 28747
rect 5994 28744 6000 28756
rect 5583 28716 6000 28744
rect 5583 28713 5595 28716
rect 5537 28707 5595 28713
rect 5994 28704 6000 28716
rect 6052 28704 6058 28756
rect 7834 28704 7840 28756
rect 7892 28744 7898 28756
rect 8205 28747 8263 28753
rect 8205 28744 8217 28747
rect 7892 28716 8217 28744
rect 7892 28704 7898 28716
rect 8205 28713 8217 28716
rect 8251 28713 8263 28747
rect 18598 28744 18604 28756
rect 18559 28716 18604 28744
rect 8205 28707 8263 28713
rect 18598 28704 18604 28716
rect 18656 28704 18662 28756
rect 26789 28747 26847 28753
rect 26789 28713 26801 28747
rect 26835 28744 26847 28747
rect 27154 28744 27160 28756
rect 26835 28716 27160 28744
rect 26835 28713 26847 28716
rect 26789 28707 26847 28713
rect 27154 28704 27160 28716
rect 27212 28704 27218 28756
rect 27430 28744 27436 28756
rect 27391 28716 27436 28744
rect 27430 28704 27436 28716
rect 27488 28704 27494 28756
rect 36265 28747 36323 28753
rect 36265 28713 36277 28747
rect 36311 28744 36323 28747
rect 37550 28744 37556 28756
rect 36311 28716 37556 28744
rect 36311 28713 36323 28716
rect 36265 28707 36323 28713
rect 37550 28704 37556 28716
rect 37608 28704 37614 28756
rect 4982 28636 4988 28688
rect 5040 28676 5046 28688
rect 5353 28679 5411 28685
rect 5353 28676 5365 28679
rect 5040 28648 5365 28676
rect 5040 28636 5046 28648
rect 5353 28645 5365 28648
rect 5399 28645 5411 28679
rect 5353 28639 5411 28645
rect 9674 28568 9680 28620
rect 9732 28608 9738 28620
rect 14277 28611 14335 28617
rect 14277 28608 14289 28611
rect 9732 28580 14289 28608
rect 9732 28568 9738 28580
rect 14277 28577 14289 28580
rect 14323 28608 14335 28611
rect 14550 28608 14556 28620
rect 14323 28580 14556 28608
rect 14323 28577 14335 28580
rect 14277 28571 14335 28577
rect 14550 28568 14556 28580
rect 14608 28568 14614 28620
rect 5077 28543 5135 28549
rect 5077 28509 5089 28543
rect 5123 28540 5135 28543
rect 5350 28540 5356 28552
rect 5123 28512 5356 28540
rect 5123 28509 5135 28512
rect 5077 28503 5135 28509
rect 5350 28500 5356 28512
rect 5408 28500 5414 28552
rect 6178 28540 6184 28552
rect 6139 28512 6184 28540
rect 6178 28500 6184 28512
rect 6236 28500 6242 28552
rect 6270 28500 6276 28552
rect 6328 28540 6334 28552
rect 6365 28543 6423 28549
rect 6365 28540 6377 28543
rect 6328 28512 6377 28540
rect 6328 28500 6334 28512
rect 6365 28509 6377 28512
rect 6411 28509 6423 28543
rect 6365 28503 6423 28509
rect 6730 28500 6736 28552
rect 6788 28540 6794 28552
rect 7006 28540 7012 28552
rect 6788 28512 7012 28540
rect 6788 28500 6794 28512
rect 7006 28500 7012 28512
rect 7064 28500 7070 28552
rect 7285 28543 7343 28549
rect 7285 28509 7297 28543
rect 7331 28509 7343 28543
rect 7926 28540 7932 28552
rect 7887 28512 7932 28540
rect 7285 28503 7343 28509
rect 4338 28432 4344 28484
rect 4396 28472 4402 28484
rect 4433 28475 4491 28481
rect 4433 28472 4445 28475
rect 4396 28444 4445 28472
rect 4396 28432 4402 28444
rect 4433 28441 4445 28444
rect 4479 28441 4491 28475
rect 7300 28472 7328 28503
rect 7926 28500 7932 28512
rect 7984 28500 7990 28552
rect 14366 28540 14372 28552
rect 14327 28512 14372 28540
rect 14366 28500 14372 28512
rect 14424 28500 14430 28552
rect 17770 28500 17776 28552
rect 17828 28540 17834 28552
rect 19245 28543 19303 28549
rect 19245 28540 19257 28543
rect 17828 28512 19257 28540
rect 17828 28500 17834 28512
rect 19245 28509 19257 28512
rect 19291 28509 19303 28543
rect 26786 28540 26792 28552
rect 26747 28512 26792 28540
rect 19245 28503 19303 28509
rect 26786 28500 26792 28512
rect 26844 28500 26850 28552
rect 27522 28540 27528 28552
rect 27483 28512 27528 28540
rect 27522 28500 27528 28512
rect 27580 28500 27586 28552
rect 35069 28543 35127 28549
rect 35069 28509 35081 28543
rect 35115 28509 35127 28543
rect 35342 28540 35348 28552
rect 35303 28512 35348 28540
rect 35069 28503 35127 28509
rect 7650 28472 7656 28484
rect 7300 28444 7656 28472
rect 4433 28435 4491 28441
rect 7650 28432 7656 28444
rect 7708 28472 7714 28484
rect 7708 28444 8892 28472
rect 7708 28432 7714 28444
rect 8864 28416 8892 28444
rect 4525 28407 4583 28413
rect 4525 28373 4537 28407
rect 4571 28404 4583 28407
rect 6454 28404 6460 28416
rect 4571 28376 6460 28404
rect 4571 28373 4583 28376
rect 4525 28367 4583 28373
rect 6454 28364 6460 28376
rect 6512 28364 6518 28416
rect 6549 28407 6607 28413
rect 6549 28373 6561 28407
rect 6595 28404 6607 28407
rect 8018 28404 8024 28416
rect 6595 28376 8024 28404
rect 6595 28373 6607 28376
rect 6549 28367 6607 28373
rect 8018 28364 8024 28376
rect 8076 28364 8082 28416
rect 8846 28364 8852 28416
rect 8904 28404 8910 28416
rect 8941 28407 8999 28413
rect 8941 28404 8953 28407
rect 8904 28376 8953 28404
rect 8904 28364 8910 28376
rect 8941 28373 8953 28376
rect 8987 28373 8999 28407
rect 9582 28404 9588 28416
rect 9543 28376 9588 28404
rect 8941 28367 8999 28373
rect 9582 28364 9588 28376
rect 9640 28364 9646 28416
rect 14737 28407 14795 28413
rect 14737 28373 14749 28407
rect 14783 28404 14795 28407
rect 15286 28404 15292 28416
rect 14783 28376 15292 28404
rect 14783 28373 14795 28376
rect 14737 28367 14795 28373
rect 15286 28364 15292 28376
rect 15344 28364 15350 28416
rect 18046 28404 18052 28416
rect 18007 28376 18052 28404
rect 18046 28364 18052 28376
rect 18104 28364 18110 28416
rect 19429 28407 19487 28413
rect 19429 28373 19441 28407
rect 19475 28404 19487 28407
rect 20346 28404 20352 28416
rect 19475 28376 20352 28404
rect 19475 28373 19487 28376
rect 19429 28367 19487 28373
rect 20346 28364 20352 28376
rect 20404 28364 20410 28416
rect 34149 28407 34207 28413
rect 34149 28373 34161 28407
rect 34195 28404 34207 28407
rect 35084 28404 35112 28503
rect 35342 28500 35348 28512
rect 35400 28500 35406 28552
rect 36081 28543 36139 28549
rect 36081 28509 36093 28543
rect 36127 28540 36139 28543
rect 36262 28540 36268 28552
rect 36127 28512 36268 28540
rect 36127 28509 36139 28512
rect 36081 28503 36139 28509
rect 36262 28500 36268 28512
rect 36320 28500 36326 28552
rect 35158 28404 35164 28416
rect 34195 28376 35164 28404
rect 34195 28373 34207 28376
rect 34149 28367 34207 28373
rect 35158 28364 35164 28376
rect 35216 28364 35222 28416
rect 1104 28314 58880 28336
rect 1104 28262 15398 28314
rect 15450 28262 15462 28314
rect 15514 28262 15526 28314
rect 15578 28262 15590 28314
rect 15642 28262 15654 28314
rect 15706 28262 29846 28314
rect 29898 28262 29910 28314
rect 29962 28262 29974 28314
rect 30026 28262 30038 28314
rect 30090 28262 30102 28314
rect 30154 28262 44294 28314
rect 44346 28262 44358 28314
rect 44410 28262 44422 28314
rect 44474 28262 44486 28314
rect 44538 28262 44550 28314
rect 44602 28262 58880 28314
rect 1104 28240 58880 28262
rect 2314 28200 2320 28212
rect 2275 28172 2320 28200
rect 2314 28160 2320 28172
rect 2372 28160 2378 28212
rect 6362 28200 6368 28212
rect 6323 28172 6368 28200
rect 6362 28160 6368 28172
rect 6420 28160 6426 28212
rect 6454 28160 6460 28212
rect 6512 28200 6518 28212
rect 18046 28200 18052 28212
rect 6512 28172 18052 28200
rect 6512 28160 6518 28172
rect 18046 28160 18052 28172
rect 18104 28200 18110 28212
rect 20622 28200 20628 28212
rect 18104 28172 20628 28200
rect 18104 28160 18110 28172
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 36357 28203 36415 28209
rect 36357 28169 36369 28203
rect 36403 28200 36415 28203
rect 37550 28200 37556 28212
rect 36403 28172 37556 28200
rect 36403 28169 36415 28172
rect 36357 28163 36415 28169
rect 37550 28160 37556 28172
rect 37608 28160 37614 28212
rect 2774 28092 2780 28144
rect 2832 28092 2838 28144
rect 3789 28135 3847 28141
rect 3789 28101 3801 28135
rect 3835 28132 3847 28135
rect 4246 28132 4252 28144
rect 3835 28104 4252 28132
rect 3835 28101 3847 28104
rect 3789 28095 3847 28101
rect 4246 28092 4252 28104
rect 4304 28092 4310 28144
rect 6270 28092 6276 28144
rect 6328 28132 6334 28144
rect 6328 28104 6914 28132
rect 6328 28092 6334 28104
rect 4985 28067 5043 28073
rect 4985 28033 4997 28067
rect 5031 28064 5043 28067
rect 5534 28064 5540 28076
rect 5031 28036 5540 28064
rect 5031 28033 5043 28036
rect 4985 28027 5043 28033
rect 5534 28024 5540 28036
rect 5592 28024 5598 28076
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28033 6791 28067
rect 6733 28027 6791 28033
rect 1854 27996 1860 28008
rect 1767 27968 1860 27996
rect 1854 27956 1860 27968
rect 1912 27996 1918 28008
rect 2498 27996 2504 28008
rect 1912 27968 2504 27996
rect 1912 27956 1918 27968
rect 2498 27956 2504 27968
rect 2556 27996 2562 28008
rect 4065 27999 4123 28005
rect 4065 27996 4077 27999
rect 2556 27968 4077 27996
rect 2556 27956 2562 27968
rect 4065 27965 4077 27968
rect 4111 27965 4123 27999
rect 6638 27996 6644 28008
rect 6599 27968 6644 27996
rect 4065 27959 4123 27965
rect 6638 27956 6644 27968
rect 6696 27956 6702 28008
rect 6748 27928 6776 28027
rect 6886 27996 6914 28104
rect 7926 28092 7932 28144
rect 7984 28132 7990 28144
rect 8205 28135 8263 28141
rect 8205 28132 8217 28135
rect 7984 28104 8217 28132
rect 7984 28092 7990 28104
rect 8205 28101 8217 28104
rect 8251 28101 8263 28135
rect 9122 28132 9128 28144
rect 9083 28104 9128 28132
rect 8205 28095 8263 28101
rect 9122 28092 9128 28104
rect 9180 28092 9186 28144
rect 18598 28092 18604 28144
rect 18656 28132 18662 28144
rect 20346 28132 20352 28144
rect 18656 28104 19182 28132
rect 20307 28104 20352 28132
rect 18656 28092 18662 28104
rect 20346 28092 20352 28104
rect 20404 28092 20410 28144
rect 7098 28024 7104 28076
rect 7156 28064 7162 28076
rect 20640 28073 20668 28160
rect 8021 28067 8079 28073
rect 8021 28064 8033 28067
rect 7156 28036 8033 28064
rect 7156 28024 7162 28036
rect 8021 28033 8033 28036
rect 8067 28033 8079 28067
rect 8021 28027 8079 28033
rect 16945 28067 17003 28073
rect 16945 28033 16957 28067
rect 16991 28064 17003 28067
rect 17865 28067 17923 28073
rect 17865 28064 17877 28067
rect 16991 28036 17877 28064
rect 16991 28033 17003 28036
rect 16945 28027 17003 28033
rect 17865 28033 17877 28036
rect 17911 28064 17923 28067
rect 20625 28067 20683 28073
rect 17911 28036 18920 28064
rect 17911 28033 17923 28036
rect 17865 28027 17923 28033
rect 9033 27999 9091 28005
rect 9033 27996 9045 27999
rect 6886 27968 9045 27996
rect 9033 27965 9045 27968
rect 9079 27965 9091 27999
rect 9033 27959 9091 27965
rect 10045 27999 10103 28005
rect 10045 27965 10057 27999
rect 10091 27996 10103 27999
rect 17770 27996 17776 28008
rect 10091 27968 12434 27996
rect 17731 27968 17776 27996
rect 10091 27965 10103 27968
rect 10045 27959 10103 27965
rect 8754 27928 8760 27940
rect 6748 27900 8760 27928
rect 8754 27888 8760 27900
rect 8812 27928 8818 27940
rect 9674 27928 9680 27940
rect 8812 27900 9680 27928
rect 8812 27888 8818 27900
rect 9674 27888 9680 27900
rect 9732 27888 9738 27940
rect 12406 27928 12434 27968
rect 17770 27956 17776 27968
rect 17828 27956 17834 28008
rect 18892 28005 18920 28036
rect 20625 28033 20637 28067
rect 20671 28033 20683 28067
rect 20625 28027 20683 28033
rect 34790 28024 34796 28076
rect 34848 28064 34854 28076
rect 35342 28064 35348 28076
rect 34848 28036 35348 28064
rect 34848 28024 34854 28036
rect 35342 28024 35348 28036
rect 35400 28064 35406 28076
rect 35437 28067 35495 28073
rect 35437 28064 35449 28067
rect 35400 28036 35449 28064
rect 35400 28024 35406 28036
rect 35437 28033 35449 28036
rect 35483 28033 35495 28067
rect 36078 28064 36084 28076
rect 36039 28036 36084 28064
rect 35437 28027 35495 28033
rect 36078 28024 36084 28036
rect 36136 28024 36142 28076
rect 58066 28064 58072 28076
rect 58027 28036 58072 28064
rect 58066 28024 58072 28036
rect 58124 28024 58130 28076
rect 18877 27999 18935 28005
rect 18877 27965 18889 27999
rect 18923 27965 18935 27999
rect 35158 27996 35164 28008
rect 35119 27968 35164 27996
rect 18877 27959 18935 27965
rect 35158 27956 35164 27968
rect 35216 27956 35222 28008
rect 18233 27931 18291 27937
rect 12406 27900 18184 27928
rect 4338 27820 4344 27872
rect 4396 27860 4402 27872
rect 4801 27863 4859 27869
rect 4801 27860 4813 27863
rect 4396 27832 4813 27860
rect 4396 27820 4402 27832
rect 4801 27829 4813 27832
rect 4847 27829 4859 27863
rect 16758 27860 16764 27872
rect 16719 27832 16764 27860
rect 4801 27823 4859 27829
rect 16758 27820 16764 27832
rect 16816 27820 16822 27872
rect 18156 27860 18184 27900
rect 18233 27897 18245 27931
rect 18279 27928 18291 27931
rect 19334 27928 19340 27940
rect 18279 27900 19340 27928
rect 18279 27897 18291 27900
rect 18233 27891 18291 27897
rect 19334 27888 19340 27900
rect 19392 27888 19398 27940
rect 57698 27888 57704 27940
rect 57756 27928 57762 27940
rect 57885 27931 57943 27937
rect 57885 27928 57897 27931
rect 57756 27900 57897 27928
rect 57756 27888 57762 27900
rect 57885 27897 57897 27900
rect 57931 27897 57943 27931
rect 57885 27891 57943 27897
rect 19610 27860 19616 27872
rect 18156 27832 19616 27860
rect 19610 27820 19616 27832
rect 19668 27820 19674 27872
rect 34701 27863 34759 27869
rect 34701 27829 34713 27863
rect 34747 27860 34759 27863
rect 34790 27860 34796 27872
rect 34747 27832 34796 27860
rect 34747 27829 34759 27832
rect 34701 27823 34759 27829
rect 34790 27820 34796 27832
rect 34848 27820 34854 27872
rect 1104 27770 58880 27792
rect 1104 27718 8174 27770
rect 8226 27718 8238 27770
rect 8290 27718 8302 27770
rect 8354 27718 8366 27770
rect 8418 27718 8430 27770
rect 8482 27718 22622 27770
rect 22674 27718 22686 27770
rect 22738 27718 22750 27770
rect 22802 27718 22814 27770
rect 22866 27718 22878 27770
rect 22930 27718 37070 27770
rect 37122 27718 37134 27770
rect 37186 27718 37198 27770
rect 37250 27718 37262 27770
rect 37314 27718 37326 27770
rect 37378 27718 51518 27770
rect 51570 27718 51582 27770
rect 51634 27718 51646 27770
rect 51698 27718 51710 27770
rect 51762 27718 51774 27770
rect 51826 27718 58880 27770
rect 1104 27696 58880 27718
rect 16012 27659 16070 27665
rect 16012 27625 16024 27659
rect 16058 27656 16070 27659
rect 16758 27656 16764 27668
rect 16058 27628 16764 27656
rect 16058 27625 16070 27628
rect 16012 27619 16070 27625
rect 16758 27616 16764 27628
rect 16816 27616 16822 27668
rect 17497 27659 17555 27665
rect 17497 27625 17509 27659
rect 17543 27656 17555 27659
rect 17770 27656 17776 27668
rect 17543 27628 17776 27656
rect 17543 27625 17555 27628
rect 17497 27619 17555 27625
rect 17770 27616 17776 27628
rect 17828 27616 17834 27668
rect 36078 27616 36084 27668
rect 36136 27656 36142 27668
rect 40954 27656 40960 27668
rect 36136 27628 40960 27656
rect 36136 27616 36142 27628
rect 40954 27616 40960 27628
rect 41012 27616 41018 27668
rect 58066 27656 58072 27668
rect 58027 27628 58072 27656
rect 58066 27616 58072 27628
rect 58124 27616 58130 27668
rect 4246 27588 4252 27600
rect 4207 27560 4252 27588
rect 4246 27548 4252 27560
rect 4304 27548 4310 27600
rect 5353 27591 5411 27597
rect 5353 27557 5365 27591
rect 5399 27588 5411 27591
rect 5399 27560 5856 27588
rect 5399 27557 5411 27560
rect 5353 27551 5411 27557
rect 2866 27480 2872 27532
rect 2924 27520 2930 27532
rect 5828 27529 5856 27560
rect 6886 27560 15884 27588
rect 5813 27523 5871 27529
rect 2924 27492 5120 27520
rect 2924 27480 2930 27492
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27452 3295 27455
rect 4246 27452 4252 27464
rect 3283 27424 4252 27452
rect 3283 27421 3295 27424
rect 3237 27415 3295 27421
rect 4246 27412 4252 27424
rect 4304 27412 4310 27464
rect 2498 27344 2504 27396
rect 2556 27344 2562 27396
rect 2961 27387 3019 27393
rect 2961 27353 2973 27387
rect 3007 27384 3019 27387
rect 3878 27384 3884 27396
rect 3007 27356 3884 27384
rect 3007 27353 3019 27356
rect 2961 27347 3019 27353
rect 3878 27344 3884 27356
rect 3936 27344 3942 27396
rect 1489 27319 1547 27325
rect 1489 27285 1501 27319
rect 1535 27316 1547 27319
rect 3694 27316 3700 27328
rect 1535 27288 3700 27316
rect 1535 27285 1547 27288
rect 1489 27279 1547 27285
rect 3694 27276 3700 27288
rect 3752 27316 3758 27328
rect 4062 27316 4068 27328
rect 3752 27288 4068 27316
rect 3752 27276 3758 27288
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 5092 27316 5120 27492
rect 5813 27489 5825 27523
rect 5859 27489 5871 27523
rect 5813 27483 5871 27489
rect 5169 27455 5227 27461
rect 5169 27421 5181 27455
rect 5215 27421 5227 27455
rect 5169 27415 5227 27421
rect 5184 27384 5212 27415
rect 5442 27412 5448 27464
rect 5500 27452 5506 27464
rect 5997 27455 6055 27461
rect 5997 27452 6009 27455
rect 5500 27424 6009 27452
rect 5500 27412 5506 27424
rect 5997 27421 6009 27424
rect 6043 27421 6055 27455
rect 5997 27415 6055 27421
rect 6886 27384 6914 27560
rect 9674 27520 9680 27532
rect 9635 27492 9680 27520
rect 9674 27480 9680 27492
rect 9732 27480 9738 27532
rect 15286 27480 15292 27532
rect 15344 27520 15350 27532
rect 15749 27523 15807 27529
rect 15749 27520 15761 27523
rect 15344 27492 15761 27520
rect 15344 27480 15350 27492
rect 15749 27489 15761 27492
rect 15795 27489 15807 27523
rect 15856 27520 15884 27560
rect 18325 27523 18383 27529
rect 18325 27520 18337 27523
rect 15856 27492 18337 27520
rect 15749 27483 15807 27489
rect 18325 27489 18337 27492
rect 18371 27489 18383 27523
rect 19610 27520 19616 27532
rect 19571 27492 19616 27520
rect 18325 27483 18383 27489
rect 19610 27480 19616 27492
rect 19668 27520 19674 27532
rect 19668 27492 22094 27520
rect 19668 27480 19674 27492
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27452 7435 27455
rect 7466 27452 7472 27464
rect 7423 27424 7472 27452
rect 7423 27421 7435 27424
rect 7377 27415 7435 27421
rect 7466 27412 7472 27424
rect 7524 27412 7530 27464
rect 7561 27455 7619 27461
rect 7561 27421 7573 27455
rect 7607 27452 7619 27455
rect 8570 27452 8576 27464
rect 7607 27424 8576 27452
rect 7607 27421 7619 27424
rect 7561 27415 7619 27421
rect 8570 27412 8576 27424
rect 8628 27412 8634 27464
rect 9398 27412 9404 27464
rect 9456 27452 9462 27464
rect 9769 27455 9827 27461
rect 9769 27452 9781 27455
rect 9456 27424 9781 27452
rect 9456 27412 9462 27424
rect 9769 27421 9781 27424
rect 9815 27452 9827 27455
rect 14366 27452 14372 27464
rect 9815 27424 14372 27452
rect 9815 27421 9827 27424
rect 9769 27415 9827 27421
rect 14366 27412 14372 27424
rect 14424 27412 14430 27464
rect 17957 27455 18015 27461
rect 17957 27421 17969 27455
rect 18003 27452 18015 27455
rect 18230 27452 18236 27464
rect 18003 27424 18236 27452
rect 18003 27421 18015 27424
rect 17957 27415 18015 27421
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 5184 27356 6914 27384
rect 7006 27344 7012 27396
rect 7064 27384 7070 27396
rect 8021 27387 8079 27393
rect 8021 27384 8033 27387
rect 7064 27356 8033 27384
rect 7064 27344 7070 27356
rect 8021 27353 8033 27356
rect 8067 27353 8079 27387
rect 8021 27347 8079 27353
rect 8205 27387 8263 27393
rect 8205 27353 8217 27387
rect 8251 27353 8263 27387
rect 8205 27347 8263 27353
rect 16408 27356 16514 27384
rect 6457 27319 6515 27325
rect 6457 27316 6469 27319
rect 5092 27288 6469 27316
rect 6457 27285 6469 27288
rect 6503 27316 6515 27319
rect 6917 27319 6975 27325
rect 6917 27316 6929 27319
rect 6503 27288 6929 27316
rect 6503 27285 6515 27288
rect 6457 27279 6515 27285
rect 6917 27285 6929 27288
rect 6963 27285 6975 27319
rect 6917 27279 6975 27285
rect 7926 27276 7932 27328
rect 7984 27316 7990 27328
rect 8220 27316 8248 27347
rect 8938 27316 8944 27328
rect 7984 27288 8248 27316
rect 8899 27288 8944 27316
rect 7984 27276 7990 27288
rect 8938 27276 8944 27288
rect 8996 27276 9002 27328
rect 9582 27276 9588 27328
rect 9640 27316 9646 27328
rect 10870 27316 10876 27328
rect 9640 27288 10876 27316
rect 9640 27276 9646 27288
rect 10870 27276 10876 27288
rect 10928 27316 10934 27328
rect 15197 27319 15255 27325
rect 15197 27316 15209 27319
rect 10928 27288 15209 27316
rect 10928 27276 10934 27288
rect 15197 27285 15209 27288
rect 15243 27316 15255 27319
rect 15746 27316 15752 27328
rect 15243 27288 15752 27316
rect 15243 27285 15255 27288
rect 15197 27279 15255 27285
rect 15746 27276 15752 27288
rect 15804 27316 15810 27328
rect 16408 27316 16436 27356
rect 18046 27344 18052 27396
rect 18104 27384 18110 27396
rect 18141 27387 18199 27393
rect 18141 27384 18153 27387
rect 18104 27356 18153 27384
rect 18104 27344 18110 27356
rect 18141 27353 18153 27356
rect 18187 27384 18199 27387
rect 19337 27387 19395 27393
rect 19337 27384 19349 27387
rect 18187 27356 19349 27384
rect 18187 27353 18199 27356
rect 18141 27347 18199 27353
rect 19337 27353 19349 27356
rect 19383 27353 19395 27387
rect 19337 27347 19395 27353
rect 19426 27344 19432 27396
rect 19484 27384 19490 27396
rect 22066 27384 22094 27492
rect 45830 27384 45836 27396
rect 19484 27356 19529 27384
rect 22066 27356 45836 27384
rect 19484 27344 19490 27356
rect 45830 27344 45836 27356
rect 45888 27344 45894 27396
rect 15804 27288 16436 27316
rect 15804 27276 15810 27288
rect 30282 27276 30288 27328
rect 30340 27316 30346 27328
rect 34977 27319 35035 27325
rect 34977 27316 34989 27319
rect 30340 27288 34989 27316
rect 30340 27276 30346 27288
rect 34977 27285 34989 27288
rect 35023 27316 35035 27319
rect 35158 27316 35164 27328
rect 35023 27288 35164 27316
rect 35023 27285 35035 27288
rect 34977 27279 35035 27285
rect 35158 27276 35164 27288
rect 35216 27276 35222 27328
rect 1104 27226 58880 27248
rect 1104 27174 15398 27226
rect 15450 27174 15462 27226
rect 15514 27174 15526 27226
rect 15578 27174 15590 27226
rect 15642 27174 15654 27226
rect 15706 27174 29846 27226
rect 29898 27174 29910 27226
rect 29962 27174 29974 27226
rect 30026 27174 30038 27226
rect 30090 27174 30102 27226
rect 30154 27174 44294 27226
rect 44346 27174 44358 27226
rect 44410 27174 44422 27226
rect 44474 27174 44486 27226
rect 44538 27174 44550 27226
rect 44602 27174 58880 27226
rect 1104 27152 58880 27174
rect 2498 27072 2504 27124
rect 2556 27112 2562 27124
rect 3237 27115 3295 27121
rect 3237 27112 3249 27115
rect 2556 27084 3249 27112
rect 2556 27072 2562 27084
rect 3237 27081 3249 27084
rect 3283 27112 3295 27115
rect 4154 27112 4160 27124
rect 3283 27084 4160 27112
rect 3283 27081 3295 27084
rect 3237 27075 3295 27081
rect 4154 27072 4160 27084
rect 4212 27072 4218 27124
rect 5442 27112 5448 27124
rect 5403 27084 5448 27112
rect 5442 27072 5448 27084
rect 5500 27072 5506 27124
rect 5534 27072 5540 27124
rect 5592 27112 5598 27124
rect 8938 27112 8944 27124
rect 5592 27084 8944 27112
rect 5592 27072 5598 27084
rect 8938 27072 8944 27084
rect 8996 27072 9002 27124
rect 18046 27112 18052 27124
rect 18007 27084 18052 27112
rect 18046 27072 18052 27084
rect 18104 27072 18110 27124
rect 3878 27044 3884 27056
rect 3839 27016 3884 27044
rect 3878 27004 3884 27016
rect 3936 27004 3942 27056
rect 4062 27004 4068 27056
rect 4120 27044 4126 27056
rect 4120 27016 5120 27044
rect 4120 27004 4126 27016
rect 3786 26936 3792 26988
rect 3844 26976 3850 26988
rect 5092 26985 5120 27016
rect 9950 27004 9956 27056
rect 10008 27044 10014 27056
rect 15105 27047 15163 27053
rect 15105 27044 15117 27047
rect 10008 27016 15117 27044
rect 10008 27004 10014 27016
rect 15105 27013 15117 27016
rect 15151 27044 15163 27047
rect 15746 27044 15752 27056
rect 15151 27016 15752 27044
rect 15151 27013 15163 27016
rect 15105 27007 15163 27013
rect 15746 27004 15752 27016
rect 15804 27004 15810 27056
rect 16853 27047 16911 27053
rect 16853 27013 16865 27047
rect 16899 27044 16911 27047
rect 17678 27044 17684 27056
rect 16899 27016 17684 27044
rect 16899 27013 16911 27016
rect 16853 27007 16911 27013
rect 17678 27004 17684 27016
rect 17736 27004 17742 27056
rect 3973 26979 4031 26985
rect 3973 26976 3985 26979
rect 3844 26948 3985 26976
rect 3844 26936 3850 26948
rect 3973 26945 3985 26948
rect 4019 26976 4031 26979
rect 5077 26979 5135 26985
rect 4019 26948 5028 26976
rect 4019 26945 4031 26948
rect 3973 26939 4031 26945
rect 5000 26917 5028 26948
rect 5077 26945 5089 26979
rect 5123 26945 5135 26979
rect 5077 26939 5135 26945
rect 7742 26936 7748 26988
rect 7800 26936 7806 26988
rect 8018 26936 8024 26988
rect 8076 26976 8082 26988
rect 8757 26979 8815 26985
rect 8757 26976 8769 26979
rect 8076 26948 8769 26976
rect 8076 26936 8082 26948
rect 8757 26945 8769 26948
rect 8803 26945 8815 26979
rect 14458 26976 14464 26988
rect 14419 26948 14464 26976
rect 8757 26939 8815 26945
rect 14458 26936 14464 26948
rect 14516 26936 14522 26988
rect 15286 26976 15292 26988
rect 15247 26948 15292 26976
rect 15286 26936 15292 26948
rect 15344 26936 15350 26988
rect 17494 26936 17500 26988
rect 17552 26976 17558 26988
rect 17865 26979 17923 26985
rect 17865 26976 17877 26979
rect 17552 26948 17877 26976
rect 17552 26936 17558 26948
rect 17865 26945 17877 26948
rect 17911 26945 17923 26979
rect 19245 26979 19303 26985
rect 19245 26976 19257 26979
rect 17865 26939 17923 26945
rect 18708 26948 19257 26976
rect 4985 26911 5043 26917
rect 4985 26877 4997 26911
rect 5031 26877 5043 26911
rect 4985 26871 5043 26877
rect 6365 26911 6423 26917
rect 6365 26877 6377 26911
rect 6411 26877 6423 26911
rect 6365 26871 6423 26877
rect 6641 26911 6699 26917
rect 6641 26877 6653 26911
rect 6687 26908 6699 26911
rect 7650 26908 7656 26920
rect 6687 26880 7656 26908
rect 6687 26877 6699 26880
rect 6641 26871 6699 26877
rect 4062 26800 4068 26852
rect 4120 26840 4126 26852
rect 6380 26840 6408 26871
rect 7650 26868 7656 26880
rect 7708 26868 7714 26920
rect 8113 26911 8171 26917
rect 8113 26877 8125 26911
rect 8159 26908 8171 26911
rect 8938 26908 8944 26920
rect 8159 26880 8944 26908
rect 8159 26877 8171 26880
rect 8113 26871 8171 26877
rect 8938 26868 8944 26880
rect 8996 26868 9002 26920
rect 14550 26908 14556 26920
rect 14511 26880 14556 26908
rect 14550 26868 14556 26880
rect 14608 26868 14614 26920
rect 15930 26868 15936 26920
rect 15988 26908 15994 26920
rect 18708 26917 18736 26948
rect 19245 26945 19257 26948
rect 19291 26945 19303 26979
rect 19245 26939 19303 26945
rect 23382 26936 23388 26988
rect 23440 26976 23446 26988
rect 23569 26979 23627 26985
rect 23569 26976 23581 26979
rect 23440 26948 23581 26976
rect 23440 26936 23446 26948
rect 23569 26945 23581 26948
rect 23615 26945 23627 26979
rect 23569 26939 23627 26945
rect 18693 26911 18751 26917
rect 18693 26908 18705 26911
rect 15988 26880 18705 26908
rect 15988 26868 15994 26880
rect 18693 26877 18705 26880
rect 18739 26877 18751 26911
rect 18693 26871 18751 26877
rect 9309 26843 9367 26849
rect 9309 26840 9321 26843
rect 4120 26812 6408 26840
rect 4120 26800 4126 26812
rect 2406 26732 2412 26784
rect 2464 26772 2470 26784
rect 2501 26775 2559 26781
rect 2501 26772 2513 26775
rect 2464 26744 2513 26772
rect 2464 26732 2470 26744
rect 2501 26741 2513 26744
rect 2547 26772 2559 26775
rect 4430 26772 4436 26784
rect 2547 26744 4436 26772
rect 2547 26741 2559 26744
rect 2501 26735 2559 26741
rect 4430 26732 4436 26744
rect 4488 26732 4494 26784
rect 6380 26772 6408 26812
rect 8036 26812 9321 26840
rect 8036 26772 8064 26812
rect 9309 26809 9321 26812
rect 9355 26840 9367 26843
rect 9858 26840 9864 26852
rect 9355 26812 9864 26840
rect 9355 26809 9367 26812
rect 9309 26803 9367 26809
rect 9858 26800 9864 26812
rect 9916 26840 9922 26852
rect 11609 26843 11667 26849
rect 11609 26840 11621 26843
rect 9916 26812 11621 26840
rect 9916 26800 9922 26812
rect 11609 26809 11621 26812
rect 11655 26840 11667 26843
rect 13633 26843 13691 26849
rect 13633 26840 13645 26843
rect 11655 26812 13645 26840
rect 11655 26809 11667 26812
rect 11609 26803 11667 26809
rect 13633 26809 13645 26812
rect 13679 26840 13691 26843
rect 13814 26840 13820 26852
rect 13679 26812 13820 26840
rect 13679 26809 13691 26812
rect 13633 26803 13691 26809
rect 13814 26800 13820 26812
rect 13872 26840 13878 26852
rect 19429 26843 19487 26849
rect 13872 26812 17448 26840
rect 13872 26800 13878 26812
rect 8570 26772 8576 26784
rect 6380 26744 8064 26772
rect 8531 26744 8576 26772
rect 8570 26732 8576 26744
rect 8628 26732 8634 26784
rect 12345 26775 12403 26781
rect 12345 26741 12357 26775
rect 12391 26772 12403 26775
rect 12526 26772 12532 26784
rect 12391 26744 12532 26772
rect 12391 26741 12403 26744
rect 12345 26735 12403 26741
rect 12526 26732 12532 26744
rect 12584 26732 12590 26784
rect 14182 26772 14188 26784
rect 14143 26744 14188 26772
rect 14182 26732 14188 26744
rect 14240 26732 14246 26784
rect 17420 26781 17448 26812
rect 19429 26809 19441 26843
rect 19475 26840 19487 26843
rect 20714 26840 20720 26852
rect 19475 26812 20720 26840
rect 19475 26809 19487 26812
rect 19429 26803 19487 26809
rect 20714 26800 20720 26812
rect 20772 26800 20778 26852
rect 23014 26800 23020 26852
rect 23072 26840 23078 26852
rect 23385 26843 23443 26849
rect 23385 26840 23397 26843
rect 23072 26812 23397 26840
rect 23072 26800 23078 26812
rect 23385 26809 23397 26812
rect 23431 26809 23443 26843
rect 23385 26803 23443 26809
rect 17405 26775 17463 26781
rect 17405 26741 17417 26775
rect 17451 26772 17463 26775
rect 17862 26772 17868 26784
rect 17451 26744 17868 26772
rect 17451 26741 17463 26744
rect 17405 26735 17463 26741
rect 17862 26732 17868 26744
rect 17920 26732 17926 26784
rect 19981 26775 20039 26781
rect 19981 26741 19993 26775
rect 20027 26772 20039 26775
rect 20070 26772 20076 26784
rect 20027 26744 20076 26772
rect 20027 26741 20039 26744
rect 19981 26735 20039 26741
rect 20070 26732 20076 26744
rect 20128 26732 20134 26784
rect 24210 26772 24216 26784
rect 24123 26744 24216 26772
rect 24210 26732 24216 26744
rect 24268 26772 24274 26784
rect 30282 26772 30288 26784
rect 24268 26744 30288 26772
rect 24268 26732 24274 26744
rect 30282 26732 30288 26744
rect 30340 26732 30346 26784
rect 1104 26682 58880 26704
rect 1104 26630 8174 26682
rect 8226 26630 8238 26682
rect 8290 26630 8302 26682
rect 8354 26630 8366 26682
rect 8418 26630 8430 26682
rect 8482 26630 22622 26682
rect 22674 26630 22686 26682
rect 22738 26630 22750 26682
rect 22802 26630 22814 26682
rect 22866 26630 22878 26682
rect 22930 26630 37070 26682
rect 37122 26630 37134 26682
rect 37186 26630 37198 26682
rect 37250 26630 37262 26682
rect 37314 26630 37326 26682
rect 37378 26630 51518 26682
rect 51570 26630 51582 26682
rect 51634 26630 51646 26682
rect 51698 26630 51710 26682
rect 51762 26630 51774 26682
rect 51826 26630 58880 26682
rect 1104 26608 58880 26630
rect 3786 26568 3792 26580
rect 3747 26540 3792 26568
rect 3786 26528 3792 26540
rect 3844 26528 3850 26580
rect 10870 26568 10876 26580
rect 10831 26540 10876 26568
rect 10870 26528 10876 26540
rect 10928 26528 10934 26580
rect 11164 26540 17172 26568
rect 5902 26460 5908 26512
rect 5960 26500 5966 26512
rect 6181 26503 6239 26509
rect 6181 26500 6193 26503
rect 5960 26472 6193 26500
rect 5960 26460 5966 26472
rect 6181 26469 6193 26472
rect 6227 26469 6239 26503
rect 6181 26463 6239 26469
rect 8018 26460 8024 26512
rect 8076 26500 8082 26512
rect 9125 26503 9183 26509
rect 9125 26500 9137 26503
rect 8076 26472 9137 26500
rect 8076 26460 8082 26472
rect 9125 26469 9137 26472
rect 9171 26500 9183 26503
rect 11164 26500 11192 26540
rect 9171 26472 11192 26500
rect 9171 26469 9183 26472
rect 9125 26463 9183 26469
rect 12250 26460 12256 26512
rect 12308 26500 12314 26512
rect 12805 26503 12863 26509
rect 12805 26500 12817 26503
rect 12308 26472 12817 26500
rect 12308 26460 12314 26472
rect 12805 26469 12817 26472
rect 12851 26469 12863 26503
rect 12805 26463 12863 26469
rect 4062 26392 4068 26444
rect 4120 26392 4126 26444
rect 5534 26432 5540 26444
rect 5495 26404 5540 26432
rect 5534 26392 5540 26404
rect 5592 26392 5598 26444
rect 5718 26392 5724 26444
rect 5776 26432 5782 26444
rect 6638 26432 6644 26444
rect 5776 26404 6644 26432
rect 5776 26392 5782 26404
rect 6638 26392 6644 26404
rect 6696 26392 6702 26444
rect 7926 26392 7932 26444
rect 7984 26432 7990 26444
rect 8113 26435 8171 26441
rect 8113 26432 8125 26435
rect 7984 26404 8125 26432
rect 7984 26392 7990 26404
rect 8113 26401 8125 26404
rect 8159 26401 8171 26435
rect 9950 26432 9956 26444
rect 8113 26395 8171 26401
rect 8404 26404 9956 26432
rect 2409 26367 2467 26373
rect 2409 26333 2421 26367
rect 2455 26364 2467 26367
rect 2866 26364 2872 26376
rect 2455 26336 2872 26364
rect 2455 26333 2467 26336
rect 2409 26327 2467 26333
rect 2866 26324 2872 26336
rect 2924 26324 2930 26376
rect 4080 26364 4108 26392
rect 5552 26364 5580 26392
rect 5810 26364 5816 26376
rect 3160 26336 4186 26364
rect 5552 26336 5816 26364
rect 1670 26188 1676 26240
rect 1728 26228 1734 26240
rect 2317 26231 2375 26237
rect 2317 26228 2329 26231
rect 1728 26200 2329 26228
rect 1728 26188 1734 26200
rect 2317 26197 2329 26200
rect 2363 26197 2375 26231
rect 2317 26191 2375 26197
rect 3050 26188 3056 26240
rect 3108 26228 3114 26240
rect 3160 26237 3188 26336
rect 5810 26324 5816 26336
rect 5868 26324 5874 26376
rect 6549 26367 6607 26373
rect 6549 26333 6561 26367
rect 6595 26364 6607 26367
rect 6595 26336 6914 26364
rect 6595 26333 6607 26336
rect 6549 26327 6607 26333
rect 5258 26296 5264 26308
rect 5219 26268 5264 26296
rect 5258 26256 5264 26268
rect 5316 26256 5322 26308
rect 6886 26296 6914 26336
rect 7742 26324 7748 26376
rect 7800 26364 7806 26376
rect 8404 26373 8432 26404
rect 9950 26392 9956 26404
rect 10008 26392 10014 26444
rect 14642 26432 14648 26444
rect 14603 26404 14648 26432
rect 14642 26392 14648 26404
rect 14700 26392 14706 26444
rect 15102 26432 15108 26444
rect 15063 26404 15108 26432
rect 15102 26392 15108 26404
rect 15160 26392 15166 26444
rect 17144 26432 17172 26540
rect 17218 26528 17224 26580
rect 17276 26568 17282 26580
rect 17497 26571 17555 26577
rect 17497 26568 17509 26571
rect 17276 26540 17509 26568
rect 17276 26528 17282 26540
rect 17497 26537 17509 26540
rect 17543 26537 17555 26571
rect 17497 26531 17555 26537
rect 17678 26528 17684 26580
rect 17736 26568 17742 26580
rect 40770 26568 40776 26580
rect 17736 26540 40776 26568
rect 17736 26528 17742 26540
rect 40770 26528 40776 26540
rect 40828 26528 40834 26580
rect 18138 26500 18144 26512
rect 18099 26472 18144 26500
rect 18138 26460 18144 26472
rect 18196 26500 18202 26512
rect 18966 26500 18972 26512
rect 18196 26472 18972 26500
rect 18196 26460 18202 26472
rect 18966 26460 18972 26472
rect 19024 26460 19030 26512
rect 23382 26460 23388 26512
rect 23440 26500 23446 26512
rect 24765 26503 24823 26509
rect 24765 26500 24777 26503
rect 23440 26472 24777 26500
rect 23440 26460 23446 26472
rect 24765 26469 24777 26472
rect 24811 26469 24823 26503
rect 24765 26463 24823 26469
rect 19521 26435 19579 26441
rect 19521 26432 19533 26435
rect 17144 26404 19533 26432
rect 19521 26401 19533 26404
rect 19567 26432 19579 26435
rect 20346 26432 20352 26444
rect 19567 26404 20352 26432
rect 19567 26401 19579 26404
rect 19521 26395 19579 26401
rect 20346 26392 20352 26404
rect 20404 26392 20410 26444
rect 22097 26435 22155 26441
rect 22097 26401 22109 26435
rect 22143 26432 22155 26435
rect 24210 26432 24216 26444
rect 22143 26404 24216 26432
rect 22143 26401 22155 26404
rect 22097 26395 22155 26401
rect 24210 26392 24216 26404
rect 24268 26392 24274 26444
rect 8389 26367 8447 26373
rect 8389 26364 8401 26367
rect 7800 26336 8401 26364
rect 7800 26324 7806 26336
rect 8389 26333 8401 26336
rect 8435 26333 8447 26367
rect 8938 26364 8944 26376
rect 8899 26336 8944 26364
rect 8389 26327 8447 26333
rect 8938 26324 8944 26336
rect 8996 26324 9002 26376
rect 9398 26364 9404 26376
rect 9140 26336 9404 26364
rect 9140 26296 9168 26336
rect 9398 26324 9404 26336
rect 9456 26324 9462 26376
rect 11054 26324 11060 26376
rect 11112 26364 11118 26376
rect 12621 26367 12679 26373
rect 12621 26364 12633 26367
rect 11112 26336 12633 26364
rect 11112 26324 11118 26336
rect 12621 26333 12633 26336
rect 12667 26333 12679 26367
rect 13354 26364 13360 26376
rect 13315 26336 13360 26364
rect 12621 26327 12679 26333
rect 13354 26324 13360 26336
rect 13412 26324 13418 26376
rect 14458 26324 14464 26376
rect 14516 26364 14522 26376
rect 14737 26367 14795 26373
rect 14737 26364 14749 26367
rect 14516 26336 14749 26364
rect 14516 26324 14522 26336
rect 14737 26333 14749 26336
rect 14783 26333 14795 26367
rect 15746 26364 15752 26376
rect 15707 26336 15752 26364
rect 14737 26327 14795 26333
rect 15746 26324 15752 26336
rect 15804 26324 15810 26376
rect 15838 26324 15844 26376
rect 15896 26364 15902 26376
rect 16577 26367 16635 26373
rect 16577 26364 16589 26367
rect 15896 26336 16589 26364
rect 15896 26324 15902 26336
rect 16577 26333 16589 26336
rect 16623 26333 16635 26367
rect 17678 26364 17684 26376
rect 17639 26336 17684 26364
rect 16577 26327 16635 26333
rect 17678 26324 17684 26336
rect 17736 26324 17742 26376
rect 19610 26364 19616 26376
rect 19571 26336 19616 26364
rect 19610 26324 19616 26336
rect 19668 26324 19674 26376
rect 20438 26364 20444 26376
rect 20399 26336 20444 26364
rect 20438 26324 20444 26336
rect 20496 26324 20502 26376
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 23506 26336 24961 26364
rect 24949 26333 24961 26336
rect 24995 26364 25007 26367
rect 27338 26364 27344 26376
rect 24995 26336 27344 26364
rect 24995 26333 25007 26336
rect 24949 26327 25007 26333
rect 27338 26324 27344 26336
rect 27396 26324 27402 26376
rect 37642 26324 37648 26376
rect 37700 26364 37706 26376
rect 38381 26367 38439 26373
rect 38381 26364 38393 26367
rect 37700 26336 38393 26364
rect 37700 26324 37706 26336
rect 38381 26333 38393 26336
rect 38427 26333 38439 26367
rect 38381 26327 38439 26333
rect 6886 26268 9168 26296
rect 9214 26256 9220 26308
rect 9272 26296 9278 26308
rect 9858 26296 9864 26308
rect 9272 26268 9864 26296
rect 9272 26256 9278 26268
rect 9858 26256 9864 26268
rect 9916 26256 9922 26308
rect 12161 26299 12219 26305
rect 12161 26265 12173 26299
rect 12207 26296 12219 26299
rect 12526 26296 12532 26308
rect 12207 26268 12532 26296
rect 12207 26265 12219 26268
rect 12161 26259 12219 26265
rect 12526 26256 12532 26268
rect 12584 26256 12590 26308
rect 13446 26296 13452 26308
rect 13407 26268 13452 26296
rect 13446 26256 13452 26268
rect 13504 26256 13510 26308
rect 15010 26256 15016 26308
rect 15068 26296 15074 26308
rect 15565 26299 15623 26305
rect 15565 26296 15577 26299
rect 15068 26268 15577 26296
rect 15068 26256 15074 26268
rect 15565 26265 15577 26268
rect 15611 26265 15623 26299
rect 22370 26296 22376 26308
rect 15565 26259 15623 26265
rect 19996 26268 22232 26296
rect 22331 26268 22376 26296
rect 3145 26231 3203 26237
rect 3145 26228 3157 26231
rect 3108 26200 3157 26228
rect 3108 26188 3114 26200
rect 3145 26197 3157 26200
rect 3191 26197 3203 26231
rect 3145 26191 3203 26197
rect 16761 26231 16819 26237
rect 16761 26197 16773 26231
rect 16807 26228 16819 26231
rect 17034 26228 17040 26240
rect 16807 26200 17040 26228
rect 16807 26197 16819 26200
rect 16761 26191 16819 26197
rect 17034 26188 17040 26200
rect 17092 26188 17098 26240
rect 19996 26237 20024 26268
rect 19981 26231 20039 26237
rect 19981 26197 19993 26231
rect 20027 26197 20039 26231
rect 20622 26228 20628 26240
rect 20583 26200 20628 26228
rect 19981 26191 20039 26197
rect 20622 26188 20628 26200
rect 20680 26188 20686 26240
rect 22204 26228 22232 26268
rect 22370 26256 22376 26268
rect 22428 26256 22434 26308
rect 37550 26256 37556 26308
rect 37608 26296 37614 26308
rect 38197 26299 38255 26305
rect 38197 26296 38209 26299
rect 37608 26268 38209 26296
rect 37608 26256 37614 26268
rect 38197 26265 38209 26268
rect 38243 26265 38255 26299
rect 38197 26259 38255 26265
rect 23106 26228 23112 26240
rect 22204 26200 23112 26228
rect 23106 26188 23112 26200
rect 23164 26188 23170 26240
rect 23842 26228 23848 26240
rect 23803 26200 23848 26228
rect 23842 26188 23848 26200
rect 23900 26188 23906 26240
rect 1104 26138 58880 26160
rect 1104 26086 15398 26138
rect 15450 26086 15462 26138
rect 15514 26086 15526 26138
rect 15578 26086 15590 26138
rect 15642 26086 15654 26138
rect 15706 26086 29846 26138
rect 29898 26086 29910 26138
rect 29962 26086 29974 26138
rect 30026 26086 30038 26138
rect 30090 26086 30102 26138
rect 30154 26086 44294 26138
rect 44346 26086 44358 26138
rect 44410 26086 44422 26138
rect 44474 26086 44486 26138
rect 44538 26086 44550 26138
rect 44602 26086 58880 26138
rect 1104 26064 58880 26086
rect 3970 25984 3976 26036
rect 4028 26024 4034 26036
rect 5169 26027 5227 26033
rect 5169 26024 5181 26027
rect 4028 25996 5181 26024
rect 4028 25984 4034 25996
rect 5169 25993 5181 25996
rect 5215 26024 5227 26027
rect 5721 26027 5779 26033
rect 5721 26024 5733 26027
rect 5215 25996 5733 26024
rect 5215 25993 5227 25996
rect 5169 25987 5227 25993
rect 5721 25993 5733 25996
rect 5767 25993 5779 26027
rect 5721 25987 5779 25993
rect 7834 25984 7840 26036
rect 7892 26024 7898 26036
rect 10965 26027 11023 26033
rect 7892 25996 10824 26024
rect 7892 25984 7898 25996
rect 1670 25956 1676 25968
rect 1631 25928 1676 25956
rect 1670 25916 1676 25928
rect 1728 25916 1734 25968
rect 9950 25916 9956 25968
rect 10008 25916 10014 25968
rect 10796 25956 10824 25996
rect 10965 25993 10977 26027
rect 11011 26024 11023 26027
rect 11054 26024 11060 26036
rect 11011 25996 11060 26024
rect 11011 25993 11023 25996
rect 10965 25987 11023 25993
rect 11054 25984 11060 25996
rect 11112 25984 11118 26036
rect 15565 26027 15623 26033
rect 15565 25993 15577 26027
rect 15611 26024 15623 26027
rect 15838 26024 15844 26036
rect 15611 25996 15844 26024
rect 15611 25993 15623 25996
rect 15565 25987 15623 25993
rect 15838 25984 15844 25996
rect 15896 25984 15902 26036
rect 19797 26027 19855 26033
rect 17972 25996 19656 26024
rect 13173 25959 13231 25965
rect 13173 25956 13185 25959
rect 10796 25928 13185 25956
rect 13173 25925 13185 25928
rect 13219 25925 13231 25959
rect 13173 25919 13231 25925
rect 14093 25959 14151 25965
rect 14093 25925 14105 25959
rect 14139 25956 14151 25959
rect 14182 25956 14188 25968
rect 14139 25928 14188 25956
rect 14139 25925 14151 25928
rect 14093 25919 14151 25925
rect 14182 25916 14188 25928
rect 14240 25916 14246 25968
rect 15378 25956 15384 25968
rect 15291 25928 15384 25956
rect 15378 25916 15384 25928
rect 15436 25956 15442 25968
rect 17972 25956 18000 25996
rect 19628 25956 19656 25996
rect 19797 25993 19809 26027
rect 19843 26024 19855 26027
rect 20438 26024 20444 26036
rect 19843 25996 20444 26024
rect 19843 25993 19855 25996
rect 19797 25987 19855 25993
rect 20438 25984 20444 25996
rect 20496 25984 20502 26036
rect 22370 26024 22376 26036
rect 22331 25996 22376 26024
rect 22370 25984 22376 25996
rect 22428 25984 22434 26036
rect 23382 25956 23388 25968
rect 15436 25928 18000 25956
rect 19550 25928 23388 25956
rect 15436 25916 15442 25928
rect 23382 25916 23388 25928
rect 23440 25916 23446 25968
rect 30282 25956 30288 25968
rect 30243 25928 30288 25956
rect 30282 25916 30288 25928
rect 30340 25916 30346 25968
rect 2774 25848 2780 25900
rect 2832 25848 2838 25900
rect 3694 25888 3700 25900
rect 3655 25860 3700 25888
rect 3694 25848 3700 25860
rect 3752 25848 3758 25900
rect 3973 25891 4031 25897
rect 3973 25857 3985 25891
rect 4019 25888 4031 25891
rect 5258 25888 5264 25900
rect 4019 25860 5264 25888
rect 4019 25857 4031 25860
rect 3973 25851 4031 25857
rect 5258 25848 5264 25860
rect 5316 25848 5322 25900
rect 5534 25848 5540 25900
rect 5592 25888 5598 25900
rect 7101 25891 7159 25897
rect 7101 25888 7113 25891
rect 5592 25860 7113 25888
rect 5592 25848 5598 25860
rect 7101 25857 7113 25860
rect 7147 25857 7159 25891
rect 7101 25851 7159 25857
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25857 7987 25891
rect 8570 25888 8576 25900
rect 8531 25860 8576 25888
rect 7929 25851 7987 25857
rect 1397 25823 1455 25829
rect 1397 25789 1409 25823
rect 1443 25789 1455 25823
rect 1397 25783 1455 25789
rect 7193 25823 7251 25829
rect 7193 25789 7205 25823
rect 7239 25820 7251 25823
rect 7374 25820 7380 25832
rect 7239 25792 7380 25820
rect 7239 25789 7251 25792
rect 7193 25783 7251 25789
rect 1412 25684 1440 25783
rect 7374 25780 7380 25792
rect 7432 25780 7438 25832
rect 2866 25712 2872 25764
rect 2924 25752 2930 25764
rect 2924 25724 3188 25752
rect 2924 25712 2930 25724
rect 3050 25684 3056 25696
rect 1412 25656 3056 25684
rect 3050 25644 3056 25656
rect 3108 25644 3114 25696
rect 3160 25693 3188 25724
rect 4798 25712 4804 25764
rect 4856 25752 4862 25764
rect 7944 25752 7972 25851
rect 8570 25848 8576 25860
rect 8628 25848 8634 25900
rect 9214 25888 9220 25900
rect 9175 25860 9220 25888
rect 9214 25848 9220 25860
rect 9272 25848 9278 25900
rect 10962 25848 10968 25900
rect 11020 25888 11026 25900
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 11020 25860 11713 25888
rect 11020 25848 11026 25860
rect 11701 25857 11713 25860
rect 11747 25857 11759 25891
rect 13814 25888 13820 25900
rect 13775 25860 13820 25888
rect 11701 25851 11759 25857
rect 13814 25848 13820 25860
rect 13872 25848 13878 25900
rect 17129 25891 17187 25897
rect 17129 25888 17141 25891
rect 15580 25860 17141 25888
rect 9493 25823 9551 25829
rect 9493 25789 9505 25823
rect 9539 25820 9551 25823
rect 10870 25820 10876 25832
rect 9539 25792 10876 25820
rect 9539 25789 9551 25792
rect 9493 25783 9551 25789
rect 10870 25780 10876 25792
rect 10928 25780 10934 25832
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 11793 25823 11851 25829
rect 11793 25820 11805 25823
rect 11112 25792 11805 25820
rect 11112 25780 11118 25792
rect 11793 25789 11805 25792
rect 11839 25820 11851 25823
rect 12250 25820 12256 25832
rect 11839 25792 12256 25820
rect 11839 25789 11851 25792
rect 11793 25783 11851 25789
rect 12250 25780 12256 25792
rect 12308 25780 12314 25832
rect 14458 25780 14464 25832
rect 14516 25820 14522 25832
rect 15580 25820 15608 25860
rect 17129 25857 17141 25860
rect 17175 25857 17187 25891
rect 17129 25851 17187 25857
rect 19610 25848 19616 25900
rect 19668 25888 19674 25900
rect 20438 25888 20444 25900
rect 19668 25860 20444 25888
rect 19668 25848 19674 25860
rect 20438 25848 20444 25860
rect 20496 25848 20502 25900
rect 22005 25891 22063 25897
rect 22005 25857 22017 25891
rect 22051 25857 22063 25891
rect 23842 25888 23848 25900
rect 23803 25860 23848 25888
rect 22005 25851 22063 25857
rect 17034 25820 17040 25832
rect 14516 25792 15608 25820
rect 16995 25792 17040 25820
rect 14516 25780 14522 25792
rect 17034 25780 17040 25792
rect 17092 25780 17098 25832
rect 17862 25780 17868 25832
rect 17920 25820 17926 25832
rect 18049 25823 18107 25829
rect 18049 25820 18061 25823
rect 17920 25792 18061 25820
rect 17920 25780 17926 25792
rect 18049 25789 18061 25792
rect 18095 25789 18107 25823
rect 18322 25820 18328 25832
rect 18283 25792 18328 25820
rect 18049 25783 18107 25789
rect 18322 25780 18328 25792
rect 18380 25780 18386 25832
rect 20346 25820 20352 25832
rect 20307 25792 20352 25820
rect 20346 25780 20352 25792
rect 20404 25780 20410 25832
rect 20898 25780 20904 25832
rect 20956 25820 20962 25832
rect 21913 25823 21971 25829
rect 21913 25820 21925 25823
rect 20956 25792 21925 25820
rect 20956 25780 20962 25792
rect 21913 25789 21925 25792
rect 21959 25789 21971 25823
rect 21913 25783 21971 25789
rect 4856 25724 7972 25752
rect 4856 25712 4862 25724
rect 12526 25712 12532 25764
rect 12584 25752 12590 25764
rect 12621 25755 12679 25761
rect 12621 25752 12633 25755
rect 12584 25724 12633 25752
rect 12584 25712 12590 25724
rect 12621 25721 12633 25724
rect 12667 25752 12679 25755
rect 13630 25752 13636 25764
rect 12667 25724 13636 25752
rect 12667 25721 12679 25724
rect 12621 25715 12679 25721
rect 13630 25712 13636 25724
rect 13688 25712 13694 25764
rect 16117 25755 16175 25761
rect 16117 25721 16129 25755
rect 16163 25752 16175 25755
rect 16666 25752 16672 25764
rect 16163 25724 16672 25752
rect 16163 25721 16175 25724
rect 16117 25715 16175 25721
rect 16666 25712 16672 25724
rect 16724 25752 16730 25764
rect 17770 25752 17776 25764
rect 16724 25724 17776 25752
rect 16724 25712 16730 25724
rect 17770 25712 17776 25724
rect 17828 25712 17834 25764
rect 20806 25752 20812 25764
rect 20767 25724 20812 25752
rect 20806 25712 20812 25724
rect 20864 25712 20870 25764
rect 21542 25712 21548 25764
rect 21600 25752 21606 25764
rect 22020 25752 22048 25851
rect 23842 25848 23848 25860
rect 23900 25848 23906 25900
rect 28629 25891 28687 25897
rect 28629 25888 28641 25891
rect 28092 25860 28641 25888
rect 23661 25755 23719 25761
rect 23661 25752 23673 25755
rect 21600 25724 23673 25752
rect 21600 25712 21606 25724
rect 23661 25721 23673 25724
rect 23707 25721 23719 25755
rect 23661 25715 23719 25721
rect 3145 25687 3203 25693
rect 3145 25653 3157 25687
rect 3191 25684 3203 25687
rect 3602 25684 3608 25696
rect 3191 25656 3608 25684
rect 3191 25653 3203 25656
rect 3145 25647 3203 25653
rect 3602 25644 3608 25656
rect 3660 25644 3666 25696
rect 3970 25644 3976 25696
rect 4028 25684 4034 25696
rect 4433 25687 4491 25693
rect 4433 25684 4445 25687
rect 4028 25656 4445 25684
rect 4028 25644 4034 25656
rect 4433 25653 4445 25656
rect 4479 25653 4491 25687
rect 6822 25684 6828 25696
rect 6783 25656 6828 25684
rect 4433 25647 4491 25653
rect 6822 25644 6828 25656
rect 6880 25644 6886 25696
rect 7282 25644 7288 25696
rect 7340 25684 7346 25696
rect 8021 25687 8079 25693
rect 8021 25684 8033 25687
rect 7340 25656 8033 25684
rect 7340 25644 7346 25656
rect 8021 25653 8033 25656
rect 8067 25653 8079 25687
rect 8662 25684 8668 25696
rect 8623 25656 8668 25684
rect 8021 25647 8079 25653
rect 8662 25644 8668 25656
rect 8720 25644 8726 25696
rect 12066 25684 12072 25696
rect 12027 25656 12072 25684
rect 12066 25644 12072 25656
rect 12124 25644 12130 25696
rect 13265 25687 13323 25693
rect 13265 25653 13277 25687
rect 13311 25684 13323 25687
rect 13538 25684 13544 25696
rect 13311 25656 13544 25684
rect 13311 25653 13323 25656
rect 13265 25647 13323 25653
rect 13538 25644 13544 25656
rect 13596 25644 13602 25696
rect 17497 25687 17555 25693
rect 17497 25653 17509 25687
rect 17543 25684 17555 25687
rect 19794 25684 19800 25696
rect 17543 25656 19800 25684
rect 17543 25653 17555 25656
rect 17497 25647 17555 25653
rect 19794 25644 19800 25656
rect 19852 25644 19858 25696
rect 27430 25644 27436 25696
rect 27488 25684 27494 25696
rect 28092 25693 28120 25860
rect 28629 25857 28641 25860
rect 28675 25857 28687 25891
rect 28629 25851 28687 25857
rect 28718 25848 28724 25900
rect 28776 25888 28782 25900
rect 31021 25891 31079 25897
rect 31021 25888 31033 25891
rect 28776 25860 31033 25888
rect 28776 25848 28782 25860
rect 31021 25857 31033 25860
rect 31067 25888 31079 25891
rect 35986 25888 35992 25900
rect 31067 25860 35992 25888
rect 31067 25857 31079 25860
rect 31021 25851 31079 25857
rect 35986 25848 35992 25860
rect 36044 25848 36050 25900
rect 28077 25687 28135 25693
rect 28077 25684 28089 25687
rect 27488 25656 28089 25684
rect 27488 25644 27494 25656
rect 28077 25653 28089 25656
rect 28123 25653 28135 25687
rect 30926 25684 30932 25696
rect 30887 25656 30932 25684
rect 28077 25647 28135 25653
rect 30926 25644 30932 25656
rect 30984 25644 30990 25696
rect 1104 25594 58880 25616
rect 1104 25542 8174 25594
rect 8226 25542 8238 25594
rect 8290 25542 8302 25594
rect 8354 25542 8366 25594
rect 8418 25542 8430 25594
rect 8482 25542 22622 25594
rect 22674 25542 22686 25594
rect 22738 25542 22750 25594
rect 22802 25542 22814 25594
rect 22866 25542 22878 25594
rect 22930 25542 37070 25594
rect 37122 25542 37134 25594
rect 37186 25542 37198 25594
rect 37250 25542 37262 25594
rect 37314 25542 37326 25594
rect 37378 25542 51518 25594
rect 51570 25542 51582 25594
rect 51634 25542 51646 25594
rect 51698 25542 51710 25594
rect 51762 25542 51774 25594
rect 51826 25542 58880 25594
rect 1104 25520 58880 25542
rect 5534 25480 5540 25492
rect 5495 25452 5540 25480
rect 5534 25440 5540 25452
rect 5592 25440 5598 25492
rect 9125 25483 9183 25489
rect 9125 25449 9137 25483
rect 9171 25480 9183 25483
rect 9398 25480 9404 25492
rect 9171 25452 9404 25480
rect 9171 25449 9183 25452
rect 9125 25443 9183 25449
rect 9398 25440 9404 25452
rect 9456 25440 9462 25492
rect 10870 25480 10876 25492
rect 10831 25452 10876 25480
rect 10870 25440 10876 25452
rect 10928 25440 10934 25492
rect 13262 25480 13268 25492
rect 12084 25452 13268 25480
rect 7193 25415 7251 25421
rect 7193 25381 7205 25415
rect 7239 25412 7251 25415
rect 9214 25412 9220 25424
rect 7239 25384 9220 25412
rect 7239 25381 7251 25384
rect 7193 25375 7251 25381
rect 9214 25372 9220 25384
rect 9272 25372 9278 25424
rect 10321 25415 10379 25421
rect 10321 25381 10333 25415
rect 10367 25412 10379 25415
rect 11146 25412 11152 25424
rect 10367 25384 11152 25412
rect 10367 25381 10379 25384
rect 10321 25375 10379 25381
rect 11146 25372 11152 25384
rect 11204 25372 11210 25424
rect 6733 25347 6791 25353
rect 6733 25313 6745 25347
rect 6779 25313 6791 25347
rect 7926 25344 7932 25356
rect 6733 25307 6791 25313
rect 6840 25316 7932 25344
rect 1673 25279 1731 25285
rect 1673 25245 1685 25279
rect 1719 25276 1731 25279
rect 2406 25276 2412 25288
rect 1719 25248 2268 25276
rect 2367 25248 2412 25276
rect 1719 25245 1731 25248
rect 1673 25239 1731 25245
rect 1486 25140 1492 25152
rect 1447 25112 1492 25140
rect 1486 25100 1492 25112
rect 1544 25100 1550 25152
rect 2240 25149 2268 25248
rect 2406 25236 2412 25248
rect 2464 25236 2470 25288
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 3160 25248 3801 25276
rect 3160 25152 3188 25248
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 4065 25211 4123 25217
rect 4065 25177 4077 25211
rect 4111 25208 4123 25211
rect 4338 25208 4344 25220
rect 4111 25180 4344 25208
rect 4111 25177 4123 25180
rect 4065 25171 4123 25177
rect 4338 25168 4344 25180
rect 4396 25168 4402 25220
rect 6748 25208 6776 25307
rect 6840 25285 6868 25316
rect 7926 25304 7932 25316
rect 7984 25304 7990 25356
rect 10045 25347 10103 25353
rect 10045 25313 10057 25347
rect 10091 25344 10103 25347
rect 11054 25344 11060 25356
rect 10091 25316 11060 25344
rect 10091 25313 10103 25316
rect 10045 25307 10103 25313
rect 11054 25304 11060 25316
rect 11112 25304 11118 25356
rect 11241 25347 11299 25353
rect 11241 25313 11253 25347
rect 11287 25344 11299 25347
rect 12084 25344 12112 25452
rect 13262 25440 13268 25452
rect 13320 25440 13326 25492
rect 16945 25483 17003 25489
rect 16945 25449 16957 25483
rect 16991 25480 17003 25483
rect 18322 25480 18328 25492
rect 16991 25452 18328 25480
rect 16991 25449 17003 25452
rect 16945 25443 17003 25449
rect 18322 25440 18328 25452
rect 18380 25440 18386 25492
rect 12158 25372 12164 25424
rect 12216 25412 12222 25424
rect 14369 25415 14427 25421
rect 14369 25412 14381 25415
rect 12216 25384 14381 25412
rect 12216 25372 12222 25384
rect 14369 25381 14381 25384
rect 14415 25381 14427 25415
rect 14369 25375 14427 25381
rect 14550 25372 14556 25424
rect 14608 25412 14614 25424
rect 14608 25384 18000 25412
rect 14608 25372 14614 25384
rect 12342 25344 12348 25356
rect 11287 25316 12112 25344
rect 12303 25316 12348 25344
rect 11287 25313 11299 25316
rect 11241 25307 11299 25313
rect 12342 25304 12348 25316
rect 12400 25304 12406 25356
rect 12618 25344 12624 25356
rect 12579 25316 12624 25344
rect 12618 25304 12624 25316
rect 12676 25304 12682 25356
rect 14844 25353 14872 25384
rect 14829 25347 14887 25353
rect 14829 25313 14841 25347
rect 14875 25313 14887 25347
rect 14829 25307 14887 25313
rect 16761 25347 16819 25353
rect 16761 25313 16773 25347
rect 16807 25344 16819 25347
rect 17586 25344 17592 25356
rect 16807 25316 17592 25344
rect 16807 25313 16819 25316
rect 16761 25307 16819 25313
rect 17586 25304 17592 25316
rect 17644 25304 17650 25356
rect 6825 25279 6883 25285
rect 6825 25245 6837 25279
rect 6871 25245 6883 25279
rect 7834 25276 7840 25288
rect 7795 25248 7840 25276
rect 6825 25239 6883 25245
rect 7834 25236 7840 25248
rect 7892 25236 7898 25288
rect 8938 25276 8944 25288
rect 8899 25248 8944 25276
rect 8938 25236 8944 25248
rect 8996 25236 9002 25288
rect 9950 25276 9956 25288
rect 9911 25248 9956 25276
rect 9950 25236 9956 25248
rect 10008 25276 10014 25288
rect 10962 25276 10968 25288
rect 10008 25248 10968 25276
rect 10008 25236 10014 25248
rect 10962 25236 10968 25248
rect 11020 25276 11026 25288
rect 11149 25279 11207 25285
rect 11149 25276 11161 25279
rect 11020 25248 11161 25276
rect 11020 25236 11026 25248
rect 11149 25245 11161 25248
rect 11195 25278 11207 25279
rect 12253 25279 12311 25285
rect 11195 25276 11284 25278
rect 12253 25276 12265 25279
rect 11195 25250 12265 25276
rect 11195 25245 11207 25250
rect 11256 25248 12265 25250
rect 11149 25239 11207 25245
rect 12253 25245 12265 25248
rect 12299 25245 12311 25279
rect 12253 25239 12311 25245
rect 13081 25279 13139 25285
rect 13081 25245 13093 25279
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 8018 25208 8024 25220
rect 4448 25180 4554 25208
rect 5920 25180 6224 25208
rect 6748 25180 8024 25208
rect 2225 25143 2283 25149
rect 2225 25109 2237 25143
rect 2271 25109 2283 25143
rect 3142 25140 3148 25152
rect 3103 25112 3148 25140
rect 2225 25103 2283 25109
rect 3142 25100 3148 25112
rect 3200 25100 3206 25152
rect 3510 25100 3516 25152
rect 3568 25140 3574 25152
rect 4448 25140 4476 25180
rect 5920 25140 5948 25180
rect 6086 25140 6092 25152
rect 3568 25112 5948 25140
rect 6047 25112 6092 25140
rect 3568 25100 3574 25112
rect 6086 25100 6092 25112
rect 6144 25100 6150 25152
rect 6196 25140 6224 25180
rect 8018 25168 8024 25180
rect 8076 25168 8082 25220
rect 12618 25168 12624 25220
rect 12676 25208 12682 25220
rect 13096 25208 13124 25239
rect 14642 25236 14648 25288
rect 14700 25276 14706 25288
rect 14737 25279 14795 25285
rect 14737 25276 14749 25279
rect 14700 25248 14749 25276
rect 14700 25236 14706 25248
rect 14737 25245 14749 25248
rect 14783 25276 14795 25279
rect 15194 25276 15200 25288
rect 14783 25248 15200 25276
rect 14783 25245 14795 25248
rect 14737 25239 14795 25245
rect 15194 25236 15200 25248
rect 15252 25236 15258 25288
rect 16022 25276 16028 25288
rect 15983 25248 16028 25276
rect 16022 25236 16028 25248
rect 16080 25236 16086 25288
rect 16669 25279 16727 25285
rect 16669 25245 16681 25279
rect 16715 25276 16727 25279
rect 17402 25276 17408 25288
rect 16715 25248 17408 25276
rect 16715 25245 16727 25248
rect 16669 25239 16727 25245
rect 17402 25236 17408 25248
rect 17460 25236 17466 25288
rect 17770 25236 17776 25288
rect 17828 25278 17834 25288
rect 17873 25279 17931 25285
rect 17873 25278 17885 25279
rect 17828 25250 17885 25278
rect 17828 25236 17834 25250
rect 17873 25245 17885 25250
rect 17919 25245 17931 25279
rect 17972 25276 18000 25384
rect 18046 25372 18052 25424
rect 18104 25412 18110 25424
rect 19797 25415 19855 25421
rect 18104 25384 18149 25412
rect 18248 25384 19748 25412
rect 18104 25372 18110 25384
rect 18248 25276 18276 25384
rect 18322 25304 18328 25356
rect 18380 25344 18386 25356
rect 19610 25344 19616 25356
rect 18380 25316 19616 25344
rect 18380 25304 18386 25316
rect 19610 25304 19616 25316
rect 19668 25304 19674 25356
rect 19720 25344 19748 25384
rect 19797 25381 19809 25415
rect 19843 25412 19855 25415
rect 22278 25412 22284 25424
rect 19843 25384 22284 25412
rect 19843 25381 19855 25384
rect 19797 25375 19855 25381
rect 22278 25372 22284 25384
rect 22336 25372 22342 25424
rect 20990 25344 20996 25356
rect 19720 25316 20996 25344
rect 20990 25304 20996 25316
rect 21048 25304 21054 25356
rect 26326 25344 26332 25356
rect 26287 25316 26332 25344
rect 26326 25304 26332 25316
rect 26384 25304 26390 25356
rect 29825 25347 29883 25353
rect 29825 25313 29837 25347
rect 29871 25344 29883 25347
rect 31849 25347 31907 25353
rect 31849 25344 31861 25347
rect 29871 25316 31861 25344
rect 29871 25313 29883 25316
rect 29825 25307 29883 25313
rect 31849 25313 31861 25316
rect 31895 25313 31907 25347
rect 31849 25307 31907 25313
rect 17972 25248 18276 25276
rect 18693 25279 18751 25285
rect 17873 25239 17931 25245
rect 18693 25245 18705 25279
rect 18739 25276 18751 25279
rect 19702 25276 19708 25288
rect 18739 25248 19708 25276
rect 18739 25245 18751 25248
rect 18693 25239 18751 25245
rect 19702 25236 19708 25248
rect 19760 25236 19766 25288
rect 20346 25276 20352 25288
rect 20307 25248 20352 25276
rect 20346 25236 20352 25248
rect 20404 25236 20410 25288
rect 20438 25236 20444 25288
rect 20496 25276 20502 25288
rect 20533 25279 20591 25285
rect 20533 25276 20545 25279
rect 20496 25248 20545 25276
rect 20496 25236 20502 25248
rect 20533 25245 20545 25248
rect 20579 25245 20591 25279
rect 20533 25239 20591 25245
rect 21450 25236 21456 25288
rect 21508 25276 21514 25288
rect 21821 25279 21879 25285
rect 21821 25276 21833 25279
rect 21508 25248 21833 25276
rect 21508 25236 21514 25248
rect 21821 25245 21833 25248
rect 21867 25245 21879 25279
rect 21821 25239 21879 25245
rect 21910 25236 21916 25288
rect 21968 25276 21974 25288
rect 22005 25279 22063 25285
rect 22005 25276 22017 25279
rect 21968 25248 22017 25276
rect 21968 25236 21974 25248
rect 22005 25245 22017 25248
rect 22051 25245 22063 25279
rect 28718 25276 28724 25288
rect 28679 25248 28724 25276
rect 22005 25239 22063 25245
rect 28718 25236 28724 25248
rect 28776 25236 28782 25288
rect 29546 25276 29552 25288
rect 29507 25248 29552 25276
rect 29546 25236 29552 25248
rect 29604 25236 29610 25288
rect 30926 25236 30932 25288
rect 30984 25236 30990 25288
rect 31754 25276 31760 25288
rect 31715 25248 31760 25276
rect 31754 25236 31760 25248
rect 31812 25236 31818 25288
rect 34974 25276 34980 25288
rect 34935 25248 34980 25276
rect 34974 25236 34980 25248
rect 35032 25236 35038 25288
rect 19429 25211 19487 25217
rect 12676 25180 16055 25208
rect 12676 25168 12682 25180
rect 7006 25140 7012 25152
rect 6196 25112 7012 25140
rect 7006 25100 7012 25112
rect 7064 25100 7070 25152
rect 8205 25143 8263 25149
rect 8205 25109 8217 25143
rect 8251 25140 8263 25143
rect 11422 25140 11428 25152
rect 8251 25112 11428 25140
rect 8251 25109 8263 25112
rect 8205 25103 8263 25109
rect 11422 25100 11428 25112
rect 11480 25100 11486 25152
rect 12894 25100 12900 25152
rect 12952 25140 12958 25152
rect 13173 25143 13231 25149
rect 13173 25140 13185 25143
rect 12952 25112 13185 25140
rect 12952 25100 12958 25112
rect 13173 25109 13185 25112
rect 13219 25109 13231 25143
rect 15930 25140 15936 25152
rect 15891 25112 15936 25140
rect 13173 25103 13231 25109
rect 15930 25100 15936 25112
rect 15988 25100 15994 25152
rect 16027 25140 16055 25180
rect 18064 25180 19380 25208
rect 18064 25140 18092 25180
rect 16027 25112 18092 25140
rect 18601 25143 18659 25149
rect 18601 25109 18613 25143
rect 18647 25140 18659 25143
rect 18690 25140 18696 25152
rect 18647 25112 18696 25140
rect 18647 25109 18659 25112
rect 18601 25103 18659 25109
rect 18690 25100 18696 25112
rect 18748 25100 18754 25152
rect 19352 25140 19380 25180
rect 19429 25177 19441 25211
rect 19475 25208 19487 25211
rect 19518 25208 19524 25220
rect 19475 25180 19524 25208
rect 19475 25177 19487 25180
rect 19429 25171 19487 25177
rect 19518 25168 19524 25180
rect 19576 25168 19582 25220
rect 19613 25211 19671 25217
rect 19613 25177 19625 25211
rect 19659 25208 19671 25211
rect 20070 25208 20076 25220
rect 19659 25180 20076 25208
rect 19659 25177 19671 25180
rect 19613 25171 19671 25177
rect 20070 25168 20076 25180
rect 20128 25208 20134 25220
rect 22189 25211 22247 25217
rect 20128 25180 22048 25208
rect 20128 25168 20134 25180
rect 22020 25152 22048 25180
rect 22189 25177 22201 25211
rect 22235 25208 22247 25211
rect 23934 25208 23940 25220
rect 22235 25180 23940 25208
rect 22235 25177 22247 25180
rect 22189 25171 22247 25177
rect 23934 25168 23940 25180
rect 23992 25168 23998 25220
rect 26602 25208 26608 25220
rect 26563 25180 26608 25208
rect 26602 25168 26608 25180
rect 26660 25168 26666 25220
rect 28629 25211 28687 25217
rect 28629 25208 28641 25211
rect 27830 25180 28641 25208
rect 28629 25177 28641 25180
rect 28675 25177 28687 25211
rect 28629 25171 28687 25177
rect 34514 25168 34520 25220
rect 34572 25208 34578 25220
rect 34701 25211 34759 25217
rect 34701 25208 34713 25211
rect 34572 25180 34713 25208
rect 34572 25168 34578 25180
rect 34701 25177 34713 25180
rect 34747 25177 34759 25211
rect 34701 25171 34759 25177
rect 21266 25140 21272 25152
rect 19352 25112 21272 25140
rect 21266 25100 21272 25112
rect 21324 25100 21330 25152
rect 21361 25143 21419 25149
rect 21361 25109 21373 25143
rect 21407 25140 21419 25143
rect 21450 25140 21456 25152
rect 21407 25112 21456 25140
rect 21407 25109 21419 25112
rect 21361 25103 21419 25109
rect 21450 25100 21456 25112
rect 21508 25100 21514 25152
rect 22002 25100 22008 25152
rect 22060 25100 22066 25152
rect 23017 25143 23075 25149
rect 23017 25109 23029 25143
rect 23063 25140 23075 25143
rect 23198 25140 23204 25152
rect 23063 25112 23204 25140
rect 23063 25109 23075 25112
rect 23017 25103 23075 25109
rect 23198 25100 23204 25112
rect 23256 25100 23262 25152
rect 28074 25140 28080 25152
rect 28035 25112 28080 25140
rect 28074 25100 28080 25112
rect 28132 25100 28138 25152
rect 31294 25140 31300 25152
rect 31255 25112 31300 25140
rect 31294 25100 31300 25112
rect 31352 25100 31358 25152
rect 1104 25050 58880 25072
rect 1104 24998 15398 25050
rect 15450 24998 15462 25050
rect 15514 24998 15526 25050
rect 15578 24998 15590 25050
rect 15642 24998 15654 25050
rect 15706 24998 29846 25050
rect 29898 24998 29910 25050
rect 29962 24998 29974 25050
rect 30026 24998 30038 25050
rect 30090 24998 30102 25050
rect 30154 24998 44294 25050
rect 44346 24998 44358 25050
rect 44410 24998 44422 25050
rect 44474 24998 44486 25050
rect 44538 24998 44550 25050
rect 44602 24998 58880 25050
rect 1104 24976 58880 24998
rect 4338 24896 4344 24948
rect 4396 24936 4402 24948
rect 5261 24939 5319 24945
rect 5261 24936 5273 24939
rect 4396 24908 5273 24936
rect 4396 24896 4402 24908
rect 5261 24905 5273 24908
rect 5307 24905 5319 24939
rect 16022 24936 16028 24948
rect 5261 24899 5319 24905
rect 14936 24908 16028 24936
rect 6086 24868 6092 24880
rect 5460 24840 6092 24868
rect 3694 24800 3700 24812
rect 3655 24772 3700 24800
rect 3694 24760 3700 24772
rect 3752 24760 3758 24812
rect 4798 24800 4804 24812
rect 4759 24772 4804 24800
rect 4798 24760 4804 24772
rect 4856 24760 4862 24812
rect 3602 24732 3608 24744
rect 3563 24704 3608 24732
rect 3602 24692 3608 24704
rect 3660 24692 3666 24744
rect 5460 24732 5488 24840
rect 6086 24828 6092 24840
rect 6144 24828 6150 24880
rect 7282 24868 7288 24880
rect 6748 24840 7288 24868
rect 5626 24800 5632 24812
rect 5587 24772 5632 24800
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 6748 24809 6776 24840
rect 7282 24828 7288 24840
rect 7340 24828 7346 24880
rect 9674 24868 9680 24880
rect 8588 24840 9680 24868
rect 6733 24803 6791 24809
rect 6733 24769 6745 24803
rect 6779 24769 6791 24803
rect 8588 24800 8616 24840
rect 9674 24828 9680 24840
rect 9732 24828 9738 24880
rect 12618 24868 12624 24880
rect 12579 24840 12624 24868
rect 12618 24828 12624 24840
rect 12676 24828 12682 24880
rect 12256 24812 12308 24818
rect 8142 24772 8616 24800
rect 6733 24763 6791 24769
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 8941 24803 8999 24809
rect 8941 24800 8953 24803
rect 8720 24772 8953 24800
rect 8720 24760 8726 24772
rect 8941 24769 8953 24772
rect 8987 24769 8999 24803
rect 8941 24763 8999 24769
rect 10962 24760 10968 24812
rect 11020 24800 11026 24812
rect 11609 24803 11667 24809
rect 11609 24800 11621 24803
rect 11020 24772 11621 24800
rect 11020 24760 11026 24772
rect 11609 24769 11621 24772
rect 11655 24769 11667 24803
rect 11609 24763 11667 24769
rect 12894 24760 12900 24812
rect 12952 24800 12958 24812
rect 13357 24803 13415 24809
rect 13357 24800 13369 24803
rect 12952 24772 13369 24800
rect 12952 24760 12958 24772
rect 13357 24769 13369 24772
rect 13403 24769 13415 24803
rect 13357 24763 13415 24769
rect 14185 24803 14243 24809
rect 14185 24769 14197 24803
rect 14231 24800 14243 24803
rect 14936 24800 14964 24908
rect 16022 24896 16028 24908
rect 16080 24896 16086 24948
rect 20901 24939 20959 24945
rect 20901 24905 20913 24939
rect 20947 24936 20959 24939
rect 21818 24936 21824 24948
rect 20947 24908 21824 24936
rect 20947 24905 20959 24908
rect 20901 24899 20959 24905
rect 21818 24896 21824 24908
rect 21876 24896 21882 24948
rect 22002 24896 22008 24948
rect 22060 24936 22066 24948
rect 22370 24936 22376 24948
rect 22060 24908 22376 24936
rect 22060 24896 22066 24908
rect 22370 24896 22376 24908
rect 22428 24896 22434 24948
rect 26329 24939 26387 24945
rect 26329 24905 26341 24939
rect 26375 24936 26387 24939
rect 26602 24936 26608 24948
rect 26375 24908 26608 24936
rect 26375 24905 26387 24908
rect 26329 24899 26387 24905
rect 26602 24896 26608 24908
rect 26660 24896 26666 24948
rect 19794 24828 19800 24880
rect 19852 24868 19858 24880
rect 29546 24868 29552 24880
rect 19852 24840 29552 24868
rect 19852 24828 19858 24840
rect 29546 24828 29552 24840
rect 29604 24828 29610 24880
rect 14231 24772 14964 24800
rect 15013 24803 15071 24809
rect 14231 24769 14243 24772
rect 14185 24763 14243 24769
rect 15013 24769 15025 24803
rect 15059 24769 15071 24803
rect 15013 24763 15071 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 17310 24800 17316 24812
rect 16163 24772 17316 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 12256 24754 12308 24760
rect 4448 24704 5488 24732
rect 5721 24735 5779 24741
rect 3050 24664 3056 24676
rect 2963 24636 3056 24664
rect 3050 24624 3056 24636
rect 3108 24664 3114 24676
rect 4448 24664 4476 24704
rect 5721 24701 5733 24735
rect 5767 24732 5779 24735
rect 7009 24735 7067 24741
rect 5767 24704 6684 24732
rect 5767 24701 5779 24704
rect 5721 24695 5779 24701
rect 3108 24636 4476 24664
rect 4709 24667 4767 24673
rect 3108 24624 3114 24636
rect 4709 24633 4721 24667
rect 4755 24664 4767 24667
rect 6546 24664 6552 24676
rect 4755 24636 6552 24664
rect 4755 24633 4767 24636
rect 4709 24627 4767 24633
rect 6546 24624 6552 24636
rect 6604 24624 6610 24676
rect 1946 24596 1952 24608
rect 1907 24568 1952 24596
rect 1946 24556 1952 24568
rect 2004 24556 2010 24608
rect 2222 24556 2228 24608
rect 2280 24596 2286 24608
rect 2409 24599 2467 24605
rect 2409 24596 2421 24599
rect 2280 24568 2421 24596
rect 2280 24556 2286 24568
rect 2409 24565 2421 24568
rect 2455 24565 2467 24599
rect 2409 24559 2467 24565
rect 4065 24599 4123 24605
rect 4065 24565 4077 24599
rect 4111 24596 4123 24599
rect 4890 24596 4896 24608
rect 4111 24568 4896 24596
rect 4111 24565 4123 24568
rect 4065 24559 4123 24565
rect 4890 24556 4896 24568
rect 4948 24556 4954 24608
rect 6656 24596 6684 24704
rect 7009 24701 7021 24735
rect 7055 24732 7067 24735
rect 8754 24732 8760 24744
rect 7055 24704 8760 24732
rect 7055 24701 7067 24704
rect 7009 24695 7067 24701
rect 8754 24692 8760 24704
rect 8812 24692 8818 24744
rect 9214 24732 9220 24744
rect 9175 24704 9220 24732
rect 9214 24692 9220 24704
rect 9272 24692 9278 24744
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24732 13599 24735
rect 13587 24704 14872 24732
rect 13587 24701 13599 24704
rect 13541 24695 13599 24701
rect 13722 24624 13728 24676
rect 13780 24664 13786 24676
rect 14645 24667 14703 24673
rect 14645 24664 14657 24667
rect 13780 24636 14657 24664
rect 13780 24624 13786 24636
rect 14645 24633 14657 24636
rect 14691 24633 14703 24667
rect 14645 24627 14703 24633
rect 7374 24596 7380 24608
rect 6656 24568 7380 24596
rect 7374 24556 7380 24568
rect 7432 24556 7438 24608
rect 8481 24599 8539 24605
rect 8481 24565 8493 24599
rect 8527 24596 8539 24599
rect 9674 24596 9680 24608
rect 8527 24568 9680 24596
rect 8527 24565 8539 24568
rect 8481 24559 8539 24565
rect 9674 24556 9680 24568
rect 9732 24556 9738 24608
rect 10686 24596 10692 24608
rect 10647 24568 10692 24596
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 14090 24596 14096 24608
rect 14051 24568 14096 24596
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14844 24596 14872 24704
rect 14918 24692 14924 24744
rect 14976 24732 14982 24744
rect 15028 24732 15056 24763
rect 17310 24760 17316 24772
rect 17368 24760 17374 24812
rect 17497 24803 17555 24809
rect 17497 24769 17509 24803
rect 17543 24800 17555 24803
rect 18322 24800 18328 24812
rect 17543 24772 18328 24800
rect 17543 24769 17555 24772
rect 17497 24763 17555 24769
rect 18322 24760 18328 24772
rect 18380 24760 18386 24812
rect 18693 24803 18751 24809
rect 18693 24769 18705 24803
rect 18739 24800 18751 24803
rect 18782 24800 18788 24812
rect 18739 24772 18788 24800
rect 18739 24769 18751 24772
rect 18693 24763 18751 24769
rect 18782 24760 18788 24772
rect 18840 24760 18846 24812
rect 18877 24803 18935 24809
rect 18877 24769 18889 24803
rect 18923 24800 18935 24803
rect 19150 24800 19156 24812
rect 18923 24772 19156 24800
rect 18923 24769 18935 24772
rect 18877 24763 18935 24769
rect 19150 24760 19156 24772
rect 19208 24760 19214 24812
rect 19521 24803 19579 24809
rect 19521 24769 19533 24803
rect 19567 24769 19579 24803
rect 19521 24763 19579 24769
rect 14976 24704 15056 24732
rect 15105 24735 15163 24741
rect 14976 24692 14982 24704
rect 15105 24701 15117 24735
rect 15151 24732 15163 24735
rect 15194 24732 15200 24744
rect 15151 24704 15200 24732
rect 15151 24701 15163 24704
rect 15105 24695 15163 24701
rect 15194 24692 15200 24704
rect 15252 24732 15258 24744
rect 17034 24732 17040 24744
rect 15252 24704 17040 24732
rect 15252 24692 15258 24704
rect 17034 24692 17040 24704
rect 17092 24692 17098 24744
rect 17586 24732 17592 24744
rect 17547 24704 17592 24732
rect 17586 24692 17592 24704
rect 17644 24692 17650 24744
rect 18340 24732 18368 24760
rect 19536 24732 19564 24763
rect 21266 24760 21272 24812
rect 21324 24800 21330 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21324 24772 21833 24800
rect 21324 24760 21330 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 22002 24800 22008 24812
rect 21963 24772 22008 24800
rect 21821 24763 21879 24769
rect 18340 24704 19564 24732
rect 19610 24692 19616 24744
rect 19668 24732 19674 24744
rect 20622 24732 20628 24744
rect 19668 24704 20628 24732
rect 19668 24692 19674 24704
rect 20622 24692 20628 24704
rect 20680 24692 20686 24744
rect 20993 24735 21051 24741
rect 20993 24701 21005 24735
rect 21039 24701 21051 24735
rect 20993 24695 21051 24701
rect 18506 24664 18512 24676
rect 15764 24636 18512 24664
rect 15764 24596 15792 24636
rect 18506 24624 18512 24636
rect 18564 24624 18570 24676
rect 18877 24667 18935 24673
rect 18877 24633 18889 24667
rect 18923 24664 18935 24667
rect 21008 24664 21036 24695
rect 21082 24692 21088 24744
rect 21140 24732 21146 24744
rect 21836 24732 21864 24763
rect 22002 24760 22008 24772
rect 22060 24800 22066 24812
rect 23753 24803 23811 24809
rect 23753 24800 23765 24803
rect 22060 24772 23765 24800
rect 22060 24760 22066 24772
rect 23753 24769 23765 24772
rect 23799 24769 23811 24803
rect 24486 24800 24492 24812
rect 24447 24772 24492 24800
rect 23753 24763 23811 24769
rect 24486 24760 24492 24772
rect 24544 24760 24550 24812
rect 25038 24760 25044 24812
rect 25096 24800 25102 24812
rect 25133 24803 25191 24809
rect 25133 24800 25145 24803
rect 25096 24772 25145 24800
rect 25096 24760 25102 24772
rect 25133 24769 25145 24772
rect 25179 24769 25191 24803
rect 26418 24800 26424 24812
rect 26379 24772 26424 24800
rect 25133 24763 25191 24769
rect 26418 24760 26424 24772
rect 26476 24760 26482 24812
rect 27433 24803 27491 24809
rect 27433 24769 27445 24803
rect 27479 24800 27491 24803
rect 28074 24800 28080 24812
rect 27479 24772 28080 24800
rect 27479 24769 27491 24772
rect 27433 24763 27491 24769
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 28445 24803 28503 24809
rect 28445 24769 28457 24803
rect 28491 24769 28503 24803
rect 28994 24800 29000 24812
rect 28955 24772 29000 24800
rect 28445 24763 28503 24769
rect 21910 24732 21916 24744
rect 21140 24704 21185 24732
rect 21823 24704 21916 24732
rect 21140 24692 21146 24704
rect 21910 24692 21916 24704
rect 21968 24732 21974 24744
rect 22465 24735 22523 24741
rect 22465 24732 22477 24735
rect 21968 24704 22477 24732
rect 21968 24692 21974 24704
rect 22465 24701 22477 24704
rect 22511 24701 22523 24735
rect 22465 24695 22523 24701
rect 22741 24735 22799 24741
rect 22741 24701 22753 24735
rect 22787 24732 22799 24735
rect 23382 24732 23388 24744
rect 22787 24704 23388 24732
rect 22787 24701 22799 24704
rect 22741 24695 22799 24701
rect 23382 24692 23388 24704
rect 23440 24692 23446 24744
rect 25314 24732 25320 24744
rect 25275 24704 25320 24732
rect 25314 24692 25320 24704
rect 25372 24692 25378 24744
rect 22186 24664 22192 24676
rect 18923 24636 20944 24664
rect 21008 24636 22192 24664
rect 18923 24633 18935 24636
rect 18877 24627 18935 24633
rect 14844 24568 15792 24596
rect 15838 24556 15844 24608
rect 15896 24596 15902 24608
rect 16025 24599 16083 24605
rect 16025 24596 16037 24599
rect 15896 24568 16037 24596
rect 15896 24556 15902 24568
rect 16025 24565 16037 24568
rect 16071 24565 16083 24599
rect 16025 24559 16083 24565
rect 16114 24556 16120 24608
rect 16172 24596 16178 24608
rect 17221 24599 17279 24605
rect 17221 24596 17233 24599
rect 16172 24568 17233 24596
rect 16172 24556 16178 24568
rect 17221 24565 17233 24568
rect 17267 24565 17279 24599
rect 18138 24596 18144 24608
rect 18099 24568 18144 24596
rect 17221 24559 17279 24565
rect 18138 24556 18144 24568
rect 18196 24556 18202 24608
rect 19886 24596 19892 24608
rect 19847 24568 19892 24596
rect 19886 24556 19892 24568
rect 19944 24556 19950 24608
rect 20530 24596 20536 24608
rect 20491 24568 20536 24596
rect 20530 24556 20536 24568
rect 20588 24556 20594 24608
rect 20916 24596 20944 24636
rect 22186 24624 22192 24636
rect 22244 24624 22250 24676
rect 28460 24664 28488 24763
rect 28994 24760 29000 24772
rect 29052 24760 29058 24812
rect 30009 24803 30067 24809
rect 30009 24769 30021 24803
rect 30055 24769 30067 24803
rect 30009 24763 30067 24769
rect 30929 24803 30987 24809
rect 30929 24769 30941 24803
rect 30975 24800 30987 24803
rect 31754 24800 31760 24812
rect 30975 24772 31760 24800
rect 30975 24769 30987 24772
rect 30929 24763 30987 24769
rect 30024 24732 30052 24763
rect 31754 24760 31760 24772
rect 31812 24760 31818 24812
rect 35897 24803 35955 24809
rect 35897 24800 35909 24803
rect 35006 24772 35909 24800
rect 35897 24769 35909 24772
rect 35943 24769 35955 24803
rect 35897 24763 35955 24769
rect 35986 24760 35992 24812
rect 36044 24800 36050 24812
rect 39022 24800 39028 24812
rect 36044 24772 36089 24800
rect 38778 24772 39028 24800
rect 36044 24760 36050 24772
rect 39022 24760 39028 24772
rect 39080 24760 39086 24812
rect 31021 24735 31079 24741
rect 31021 24732 31033 24735
rect 30024 24704 31033 24732
rect 31021 24701 31033 24704
rect 31067 24732 31079 24735
rect 31294 24732 31300 24744
rect 31067 24704 31300 24732
rect 31067 24701 31079 24704
rect 31021 24695 31079 24701
rect 31294 24692 31300 24704
rect 31352 24692 31358 24744
rect 31573 24735 31631 24741
rect 31573 24701 31585 24735
rect 31619 24732 31631 24735
rect 33410 24732 33416 24744
rect 31619 24704 33416 24732
rect 31619 24701 31631 24704
rect 31573 24695 31631 24701
rect 33410 24692 33416 24704
rect 33468 24692 33474 24744
rect 33594 24732 33600 24744
rect 33555 24704 33600 24732
rect 33594 24692 33600 24704
rect 33652 24692 33658 24744
rect 33873 24735 33931 24741
rect 33873 24701 33885 24735
rect 33919 24732 33931 24735
rect 34514 24732 34520 24744
rect 33919 24704 34520 24732
rect 33919 24701 33931 24704
rect 33873 24695 33931 24701
rect 34514 24692 34520 24704
rect 34572 24692 34578 24744
rect 37366 24732 37372 24744
rect 37327 24704 37372 24732
rect 37366 24692 37372 24704
rect 37424 24692 37430 24744
rect 37645 24735 37703 24741
rect 37645 24701 37657 24735
rect 37691 24732 37703 24735
rect 39942 24732 39948 24744
rect 37691 24704 39948 24732
rect 37691 24701 37703 24704
rect 37645 24695 37703 24701
rect 39942 24692 39948 24704
rect 40000 24692 40006 24744
rect 31846 24664 31852 24676
rect 28460 24636 31852 24664
rect 31846 24624 31852 24636
rect 31904 24624 31910 24676
rect 21634 24596 21640 24608
rect 20916 24568 21640 24596
rect 21634 24556 21640 24568
rect 21692 24556 21698 24608
rect 21910 24596 21916 24608
rect 21871 24568 21916 24596
rect 21910 24556 21916 24568
rect 21968 24596 21974 24608
rect 23750 24596 23756 24608
rect 21968 24568 23756 24596
rect 21968 24556 21974 24568
rect 23750 24556 23756 24568
rect 23808 24556 23814 24608
rect 23842 24556 23848 24608
rect 23900 24596 23906 24608
rect 23900 24568 23945 24596
rect 23900 24556 23906 24568
rect 26786 24556 26792 24608
rect 26844 24596 26850 24608
rect 27249 24599 27307 24605
rect 27249 24596 27261 24599
rect 26844 24568 27261 24596
rect 26844 24556 26850 24568
rect 27249 24565 27261 24568
rect 27295 24565 27307 24599
rect 28350 24596 28356 24608
rect 28311 24568 28356 24596
rect 27249 24559 27307 24565
rect 28350 24556 28356 24568
rect 28408 24556 28414 24608
rect 29181 24599 29239 24605
rect 29181 24565 29193 24599
rect 29227 24596 29239 24599
rect 29730 24596 29736 24608
rect 29227 24568 29736 24596
rect 29227 24565 29239 24568
rect 29181 24559 29239 24565
rect 29730 24556 29736 24568
rect 29788 24556 29794 24608
rect 30006 24596 30012 24608
rect 29967 24568 30012 24596
rect 30006 24556 30012 24568
rect 30064 24556 30070 24608
rect 35342 24596 35348 24608
rect 35303 24568 35348 24596
rect 35342 24556 35348 24568
rect 35400 24556 35406 24608
rect 39114 24596 39120 24608
rect 39075 24568 39120 24596
rect 39114 24556 39120 24568
rect 39172 24556 39178 24608
rect 1104 24506 58880 24528
rect 1104 24454 8174 24506
rect 8226 24454 8238 24506
rect 8290 24454 8302 24506
rect 8354 24454 8366 24506
rect 8418 24454 8430 24506
rect 8482 24454 22622 24506
rect 22674 24454 22686 24506
rect 22738 24454 22750 24506
rect 22802 24454 22814 24506
rect 22866 24454 22878 24506
rect 22930 24454 37070 24506
rect 37122 24454 37134 24506
rect 37186 24454 37198 24506
rect 37250 24454 37262 24506
rect 37314 24454 37326 24506
rect 37378 24454 51518 24506
rect 51570 24454 51582 24506
rect 51634 24454 51646 24506
rect 51698 24454 51710 24506
rect 51762 24454 51774 24506
rect 51826 24454 58880 24506
rect 1104 24432 58880 24454
rect 7193 24395 7251 24401
rect 7193 24361 7205 24395
rect 7239 24392 7251 24395
rect 9861 24395 9919 24401
rect 7239 24364 8708 24392
rect 7239 24361 7251 24364
rect 7193 24355 7251 24361
rect 4801 24327 4859 24333
rect 4801 24293 4813 24327
rect 4847 24324 4859 24327
rect 5718 24324 5724 24336
rect 4847 24296 5724 24324
rect 4847 24293 4859 24296
rect 4801 24287 4859 24293
rect 4154 24256 4160 24268
rect 3804 24228 4160 24256
rect 3142 24148 3148 24200
rect 3200 24188 3206 24200
rect 3804 24197 3832 24228
rect 4154 24216 4160 24228
rect 4212 24216 4218 24268
rect 3789 24191 3847 24197
rect 3200 24160 3245 24188
rect 3200 24148 3206 24160
rect 3789 24157 3801 24191
rect 3835 24157 3847 24191
rect 3789 24151 3847 24157
rect 3973 24191 4031 24197
rect 3973 24157 3985 24191
rect 4019 24188 4031 24191
rect 4816 24188 4844 24287
rect 5718 24284 5724 24296
rect 5776 24284 5782 24336
rect 7650 24324 7656 24336
rect 7611 24296 7656 24324
rect 7650 24284 7656 24296
rect 7708 24284 7714 24336
rect 8110 24256 8116 24268
rect 8071 24228 8116 24256
rect 8110 24216 8116 24228
rect 8168 24216 8174 24268
rect 8680 24256 8708 24364
rect 9861 24361 9873 24395
rect 9907 24392 9919 24395
rect 9950 24392 9956 24404
rect 9907 24364 9956 24392
rect 9907 24361 9919 24364
rect 9861 24355 9919 24361
rect 9950 24352 9956 24364
rect 10008 24352 10014 24404
rect 10873 24395 10931 24401
rect 10873 24361 10885 24395
rect 10919 24392 10931 24395
rect 11698 24392 11704 24404
rect 10919 24364 11704 24392
rect 10919 24361 10931 24364
rect 10873 24355 10931 24361
rect 11698 24352 11704 24364
rect 11756 24392 11762 24404
rect 13354 24392 13360 24404
rect 11756 24364 13360 24392
rect 11756 24352 11762 24364
rect 13354 24352 13360 24364
rect 13412 24352 13418 24404
rect 14458 24352 14464 24404
rect 14516 24392 14522 24404
rect 14918 24392 14924 24404
rect 14516 24364 14924 24392
rect 14516 24352 14522 24364
rect 14918 24352 14924 24364
rect 14976 24392 14982 24404
rect 15473 24395 15531 24401
rect 15473 24392 15485 24395
rect 14976 24364 15485 24392
rect 14976 24352 14982 24364
rect 15473 24361 15485 24364
rect 15519 24361 15531 24395
rect 15473 24355 15531 24361
rect 8754 24284 8760 24336
rect 8812 24324 8818 24336
rect 12621 24327 12679 24333
rect 12621 24324 12633 24327
rect 8812 24296 12633 24324
rect 8812 24284 8818 24296
rect 12621 24293 12633 24296
rect 12667 24293 12679 24327
rect 12621 24287 12679 24293
rect 10686 24256 10692 24268
rect 8680 24228 9168 24256
rect 5534 24188 5540 24200
rect 4019 24160 4844 24188
rect 5495 24160 5540 24188
rect 4019 24157 4031 24160
rect 3973 24151 4031 24157
rect 2866 24120 2872 24132
rect 2438 24092 2728 24120
rect 2827 24092 2872 24120
rect 1397 24055 1455 24061
rect 1397 24021 1409 24055
rect 1443 24052 1455 24055
rect 2038 24052 2044 24064
rect 1443 24024 2044 24052
rect 1443 24021 1455 24024
rect 1397 24015 1455 24021
rect 2038 24012 2044 24024
rect 2096 24012 2102 24064
rect 2700 24052 2728 24092
rect 2866 24080 2872 24092
rect 2924 24080 2930 24132
rect 3326 24080 3332 24132
rect 3384 24120 3390 24132
rect 3988 24120 4016 24151
rect 5534 24148 5540 24160
rect 5592 24148 5598 24200
rect 5626 24148 5632 24200
rect 5684 24188 5690 24200
rect 6273 24191 6331 24197
rect 6273 24188 6285 24191
rect 5684 24160 6285 24188
rect 5684 24148 5690 24160
rect 6273 24157 6285 24160
rect 6319 24188 6331 24191
rect 7558 24188 7564 24200
rect 6319 24160 7564 24188
rect 6319 24157 6331 24160
rect 6273 24151 6331 24157
rect 7558 24148 7564 24160
rect 7616 24148 7622 24200
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 8021 24191 8079 24197
rect 8021 24188 8033 24191
rect 7892 24160 8033 24188
rect 7892 24148 7898 24160
rect 8021 24157 8033 24160
rect 8067 24188 8079 24191
rect 8067 24160 9076 24188
rect 8067 24157 8079 24160
rect 8021 24151 8079 24157
rect 3384 24092 4016 24120
rect 4617 24123 4675 24129
rect 3384 24080 3390 24092
rect 4617 24089 4629 24123
rect 4663 24120 4675 24123
rect 4890 24120 4896 24132
rect 4663 24092 4896 24120
rect 4663 24089 4675 24092
rect 4617 24083 4675 24089
rect 4890 24080 4896 24092
rect 4948 24080 4954 24132
rect 2774 24052 2780 24064
rect 2687 24024 2780 24052
rect 2774 24012 2780 24024
rect 2832 24052 2838 24064
rect 3510 24052 3516 24064
rect 2832 24024 3516 24052
rect 2832 24012 2838 24024
rect 3510 24012 3516 24024
rect 3568 24012 3574 24064
rect 3786 24052 3792 24064
rect 3747 24024 3792 24052
rect 3786 24012 3792 24024
rect 3844 24012 3850 24064
rect 9048 24061 9076 24160
rect 9140 24120 9168 24228
rect 9232 24228 10692 24256
rect 9232 24197 9260 24228
rect 10686 24216 10692 24228
rect 10744 24216 10750 24268
rect 13081 24259 13139 24265
rect 13081 24225 13093 24259
rect 13127 24256 13139 24259
rect 13262 24256 13268 24268
rect 13127 24228 13268 24256
rect 13127 24225 13139 24228
rect 13081 24219 13139 24225
rect 13262 24216 13268 24228
rect 13320 24216 13326 24268
rect 13354 24216 13360 24268
rect 13412 24256 13418 24268
rect 14277 24259 14335 24265
rect 14277 24256 14289 24259
rect 13412 24228 14289 24256
rect 13412 24216 13418 24228
rect 14277 24225 14289 24228
rect 14323 24225 14335 24259
rect 14277 24219 14335 24225
rect 14737 24259 14795 24265
rect 14737 24225 14749 24259
rect 14783 24256 14795 24259
rect 14783 24228 15424 24256
rect 14783 24225 14795 24228
rect 14737 24219 14795 24225
rect 9217 24191 9275 24197
rect 9217 24157 9229 24191
rect 9263 24157 9275 24191
rect 9674 24188 9680 24200
rect 9635 24160 9680 24188
rect 9217 24151 9275 24157
rect 9674 24148 9680 24160
rect 9732 24148 9738 24200
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 12989 24191 13047 24197
rect 12989 24188 13001 24191
rect 12308 24160 13001 24188
rect 12308 24148 12314 24160
rect 12989 24157 13001 24160
rect 13035 24157 13047 24191
rect 14642 24188 14648 24200
rect 14603 24160 14648 24188
rect 12989 24151 13047 24157
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 15286 24188 15292 24200
rect 15247 24160 15292 24188
rect 15286 24148 15292 24160
rect 15344 24148 15350 24200
rect 10962 24120 10968 24132
rect 9140 24092 10968 24120
rect 10962 24080 10968 24092
rect 11020 24080 11026 24132
rect 12161 24123 12219 24129
rect 12161 24089 12173 24123
rect 12207 24120 12219 24123
rect 15194 24120 15200 24132
rect 12207 24092 15200 24120
rect 12207 24089 12219 24092
rect 12161 24083 12219 24089
rect 15194 24080 15200 24092
rect 15252 24080 15258 24132
rect 15396 24120 15424 24228
rect 15488 24188 15516 24355
rect 17586 24352 17592 24404
rect 17644 24392 17650 24404
rect 23293 24395 23351 24401
rect 23293 24392 23305 24395
rect 17644 24364 23305 24392
rect 17644 24352 17650 24364
rect 23293 24361 23305 24364
rect 23339 24361 23351 24395
rect 23293 24355 23351 24361
rect 23382 24352 23388 24404
rect 23440 24392 23446 24404
rect 23477 24395 23535 24401
rect 23477 24392 23489 24395
rect 23440 24364 23489 24392
rect 23440 24352 23446 24364
rect 23477 24361 23489 24364
rect 23523 24361 23535 24395
rect 25685 24395 25743 24401
rect 25685 24392 25697 24395
rect 23477 24355 23535 24361
rect 23584 24364 25697 24392
rect 22002 24324 22008 24336
rect 17328 24296 22008 24324
rect 17328 24265 17356 24296
rect 22002 24284 22008 24296
rect 22060 24284 22066 24336
rect 23584 24324 23612 24364
rect 25685 24361 25697 24364
rect 25731 24361 25743 24395
rect 25685 24355 25743 24361
rect 25130 24324 25136 24336
rect 22204 24296 23612 24324
rect 23676 24296 25136 24324
rect 17313 24259 17371 24265
rect 17313 24225 17325 24259
rect 17359 24225 17371 24259
rect 18233 24259 18291 24265
rect 18233 24256 18245 24259
rect 17313 24219 17371 24225
rect 17420 24228 18245 24256
rect 16301 24191 16359 24197
rect 16301 24188 16313 24191
rect 15488 24160 16313 24188
rect 16301 24157 16313 24160
rect 16347 24157 16359 24191
rect 17034 24188 17040 24200
rect 16974 24160 17040 24188
rect 16301 24151 16359 24157
rect 17034 24148 17040 24160
rect 17092 24148 17098 24200
rect 17420 24120 17448 24228
rect 18233 24225 18245 24228
rect 18279 24256 18291 24259
rect 18693 24259 18751 24265
rect 18279 24228 18460 24256
rect 18279 24225 18291 24228
rect 18233 24219 18291 24225
rect 18322 24188 18328 24200
rect 18283 24160 18328 24188
rect 18322 24148 18328 24160
rect 18380 24148 18386 24200
rect 18432 24188 18460 24228
rect 18693 24225 18705 24259
rect 18739 24256 18751 24259
rect 19058 24256 19064 24268
rect 18739 24228 19064 24256
rect 18739 24225 18751 24228
rect 18693 24219 18751 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 19610 24216 19616 24268
rect 19668 24216 19674 24268
rect 21818 24216 21824 24268
rect 21876 24256 21882 24268
rect 22204 24256 22232 24296
rect 21876 24228 22232 24256
rect 21876 24216 21882 24228
rect 22278 24216 22284 24268
rect 22336 24256 22342 24268
rect 22649 24259 22707 24265
rect 22649 24256 22661 24259
rect 22336 24228 22661 24256
rect 22336 24216 22342 24228
rect 22649 24225 22661 24228
rect 22695 24256 22707 24259
rect 23569 24259 23627 24265
rect 23569 24256 23581 24259
rect 22695 24228 23581 24256
rect 22695 24225 22707 24228
rect 22649 24219 22707 24225
rect 23569 24225 23581 24228
rect 23615 24225 23627 24259
rect 23569 24219 23627 24225
rect 19628 24188 19656 24216
rect 21358 24188 21364 24200
rect 18432 24160 19656 24188
rect 21319 24160 21364 24188
rect 21358 24148 21364 24160
rect 21416 24148 21422 24200
rect 22094 24148 22100 24200
rect 22152 24188 22158 24200
rect 22557 24191 22615 24197
rect 22557 24188 22569 24191
rect 22152 24160 22569 24188
rect 22152 24148 22158 24160
rect 22557 24157 22569 24160
rect 22603 24188 22615 24191
rect 23198 24188 23204 24200
rect 22603 24160 23204 24188
rect 22603 24157 22615 24160
rect 22557 24151 22615 24157
rect 23198 24148 23204 24160
rect 23256 24188 23262 24200
rect 23676 24197 23704 24296
rect 25130 24284 25136 24296
rect 25188 24284 25194 24336
rect 25700 24324 25728 24355
rect 26418 24352 26424 24404
rect 26476 24392 26482 24404
rect 27982 24392 27988 24404
rect 26476 24364 27988 24392
rect 26476 24352 26482 24364
rect 27982 24352 27988 24364
rect 28040 24392 28046 24404
rect 28261 24395 28319 24401
rect 28261 24392 28273 24395
rect 28040 24364 28273 24392
rect 28040 24352 28046 24364
rect 28261 24361 28273 24364
rect 28307 24361 28319 24395
rect 28994 24392 29000 24404
rect 28955 24364 29000 24392
rect 28261 24355 28319 24361
rect 28994 24352 29000 24364
rect 29052 24352 29058 24404
rect 30006 24352 30012 24404
rect 30064 24352 30070 24404
rect 31665 24395 31723 24401
rect 31665 24361 31677 24395
rect 31711 24392 31723 24395
rect 31754 24392 31760 24404
rect 31711 24364 31760 24392
rect 31711 24361 31723 24364
rect 31665 24355 31723 24361
rect 31754 24352 31760 24364
rect 31812 24352 31818 24404
rect 33410 24352 33416 24404
rect 33468 24392 33474 24404
rect 34149 24395 34207 24401
rect 33468 24364 33732 24392
rect 33468 24352 33474 24364
rect 25700 24296 26648 24324
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 25777 24259 25835 24265
rect 25777 24256 25789 24259
rect 24176 24228 25789 24256
rect 24176 24216 24182 24228
rect 25777 24225 25789 24228
rect 25823 24256 25835 24259
rect 26418 24256 26424 24268
rect 25823 24228 26424 24256
rect 25823 24225 25835 24228
rect 25777 24219 25835 24225
rect 26418 24216 26424 24228
rect 26476 24216 26482 24268
rect 26620 24256 26648 24296
rect 28718 24256 28724 24268
rect 26620 24228 28724 24256
rect 28718 24216 28724 24228
rect 28776 24216 28782 24268
rect 29012 24256 29040 24352
rect 29917 24259 29975 24265
rect 29917 24256 29929 24259
rect 29012 24228 29929 24256
rect 29917 24225 29929 24228
rect 29963 24225 29975 24259
rect 30024 24256 30052 24352
rect 33704 24324 33732 24364
rect 34149 24361 34161 24395
rect 34195 24392 34207 24395
rect 34974 24392 34980 24404
rect 34195 24364 34980 24392
rect 34195 24361 34207 24364
rect 34149 24355 34207 24361
rect 34974 24352 34980 24364
rect 35032 24352 35038 24404
rect 35986 24352 35992 24404
rect 36044 24392 36050 24404
rect 37734 24392 37740 24404
rect 36044 24364 37740 24392
rect 36044 24352 36050 24364
rect 37734 24352 37740 24364
rect 37792 24392 37798 24404
rect 38562 24392 38568 24404
rect 37792 24364 38568 24392
rect 37792 24352 37798 24364
rect 38562 24352 38568 24364
rect 38620 24352 38626 24404
rect 39022 24392 39028 24404
rect 38983 24364 39028 24392
rect 39022 24352 39028 24364
rect 39080 24352 39086 24404
rect 39942 24392 39948 24404
rect 39903 24364 39948 24392
rect 39942 24352 39948 24364
rect 40000 24352 40006 24404
rect 40678 24324 40684 24336
rect 33704 24296 40684 24324
rect 40678 24284 40684 24296
rect 40736 24284 40742 24336
rect 30193 24259 30251 24265
rect 30193 24256 30205 24259
rect 30024 24228 30205 24256
rect 29917 24219 29975 24225
rect 30193 24225 30205 24228
rect 30239 24225 30251 24259
rect 30193 24219 30251 24225
rect 32677 24259 32735 24265
rect 32677 24225 32689 24259
rect 32723 24256 32735 24259
rect 36541 24259 36599 24265
rect 36541 24256 36553 24259
rect 32723 24228 36553 24256
rect 32723 24225 32735 24228
rect 32677 24219 32735 24225
rect 36541 24225 36553 24228
rect 36587 24225 36599 24259
rect 39114 24256 39120 24268
rect 36541 24219 36599 24225
rect 38488 24228 39120 24256
rect 23661 24191 23719 24197
rect 23661 24188 23673 24191
rect 23256 24160 23673 24188
rect 23256 24148 23262 24160
rect 23661 24157 23673 24160
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 23750 24148 23756 24200
rect 23808 24188 23814 24200
rect 25685 24191 25743 24197
rect 25685 24188 25697 24191
rect 23808 24160 25697 24188
rect 23808 24148 23814 24160
rect 25685 24157 25697 24160
rect 25731 24157 25743 24191
rect 26510 24188 26516 24200
rect 26471 24160 26516 24188
rect 25685 24151 25743 24157
rect 26510 24148 26516 24160
rect 26568 24148 26574 24200
rect 28813 24191 28871 24197
rect 28813 24157 28825 24191
rect 28859 24188 28871 24191
rect 29546 24188 29552 24200
rect 28859 24160 29552 24188
rect 28859 24157 28871 24160
rect 28813 24151 28871 24157
rect 15396 24092 17448 24120
rect 18138 24080 18144 24132
rect 18196 24120 18202 24132
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 18196 24092 19625 24120
rect 18196 24080 18202 24092
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 19613 24083 19671 24089
rect 23842 24080 23848 24132
rect 23900 24120 23906 24132
rect 26786 24120 26792 24132
rect 23900 24092 26372 24120
rect 26747 24092 26792 24120
rect 23900 24080 23906 24092
rect 9033 24055 9091 24061
rect 9033 24021 9045 24055
rect 9079 24052 9091 24055
rect 20438 24052 20444 24064
rect 9079 24024 20444 24052
rect 9079 24021 9091 24024
rect 9033 24015 9091 24021
rect 20438 24012 20444 24024
rect 20496 24012 20502 24064
rect 20990 24012 20996 24064
rect 21048 24052 21054 24064
rect 22097 24055 22155 24061
rect 22097 24052 22109 24055
rect 21048 24024 22109 24052
rect 21048 24012 21054 24024
rect 22097 24021 22109 24024
rect 22143 24021 22155 24055
rect 22462 24052 22468 24064
rect 22423 24024 22468 24052
rect 22097 24015 22155 24021
rect 22462 24012 22468 24024
rect 22520 24012 22526 24064
rect 24489 24055 24547 24061
rect 24489 24021 24501 24055
rect 24535 24052 24547 24055
rect 24762 24052 24768 24064
rect 24535 24024 24768 24052
rect 24535 24021 24547 24024
rect 24489 24015 24547 24021
rect 24762 24012 24768 24024
rect 24820 24012 24826 24064
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 25130 24052 25136 24064
rect 25087 24024 25136 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 25130 24012 25136 24024
rect 25188 24012 25194 24064
rect 26053 24055 26111 24061
rect 26053 24021 26065 24055
rect 26099 24052 26111 24055
rect 26234 24052 26240 24064
rect 26099 24024 26240 24052
rect 26099 24021 26111 24024
rect 26053 24015 26111 24021
rect 26234 24012 26240 24024
rect 26292 24012 26298 24064
rect 26344 24052 26372 24092
rect 26786 24080 26792 24092
rect 26844 24080 26850 24132
rect 28350 24120 28356 24132
rect 28014 24092 28356 24120
rect 28350 24080 28356 24092
rect 28408 24080 28414 24132
rect 28828 24052 28856 24151
rect 29546 24148 29552 24160
rect 29604 24148 29610 24200
rect 32401 24191 32459 24197
rect 32401 24157 32413 24191
rect 32447 24157 32459 24191
rect 32401 24151 32459 24157
rect 31202 24080 31208 24132
rect 31260 24080 31266 24132
rect 26344 24024 28856 24052
rect 29454 24012 29460 24064
rect 29512 24052 29518 24064
rect 31754 24052 31760 24064
rect 29512 24024 31760 24052
rect 29512 24012 29518 24024
rect 31754 24012 31760 24024
rect 31812 24052 31818 24064
rect 32416 24052 32444 24151
rect 34974 24148 34980 24200
rect 35032 24188 35038 24200
rect 35161 24191 35219 24197
rect 35161 24188 35173 24191
rect 35032 24160 35173 24188
rect 35032 24148 35038 24160
rect 35161 24157 35173 24160
rect 35207 24157 35219 24191
rect 35161 24151 35219 24157
rect 35342 24148 35348 24200
rect 35400 24188 35406 24200
rect 38488 24197 38516 24228
rect 39114 24216 39120 24228
rect 39172 24216 39178 24268
rect 35621 24191 35679 24197
rect 35621 24188 35633 24191
rect 35400 24160 35633 24188
rect 35400 24148 35406 24160
rect 35621 24157 35633 24160
rect 35667 24188 35679 24191
rect 36449 24191 36507 24197
rect 36449 24188 36461 24191
rect 35667 24160 36461 24188
rect 35667 24157 35679 24160
rect 35621 24151 35679 24157
rect 36449 24157 36461 24160
rect 36495 24157 36507 24191
rect 36449 24151 36507 24157
rect 38473 24191 38531 24197
rect 38473 24157 38485 24191
rect 38519 24157 38531 24191
rect 38473 24151 38531 24157
rect 38562 24148 38568 24200
rect 38620 24188 38626 24200
rect 38933 24191 38991 24197
rect 38933 24188 38945 24191
rect 38620 24160 38945 24188
rect 38620 24148 38626 24160
rect 38933 24157 38945 24160
rect 38979 24157 38991 24191
rect 39850 24188 39856 24200
rect 39811 24160 39856 24188
rect 38933 24151 38991 24157
rect 39850 24148 39856 24160
rect 39908 24148 39914 24200
rect 33962 24120 33968 24132
rect 33902 24092 33968 24120
rect 33962 24080 33968 24092
rect 34020 24080 34026 24132
rect 35989 24123 36047 24129
rect 35989 24089 36001 24123
rect 36035 24120 36047 24123
rect 48314 24120 48320 24132
rect 36035 24092 48320 24120
rect 36035 24089 36047 24092
rect 35989 24083 36047 24089
rect 48314 24080 48320 24092
rect 48372 24080 48378 24132
rect 31812 24024 32444 24052
rect 31812 24012 31818 24024
rect 37550 24012 37556 24064
rect 37608 24052 37614 24064
rect 38381 24055 38439 24061
rect 38381 24052 38393 24055
rect 37608 24024 38393 24052
rect 37608 24012 37614 24024
rect 38381 24021 38393 24024
rect 38427 24021 38439 24055
rect 47578 24052 47584 24064
rect 47539 24024 47584 24052
rect 38381 24015 38439 24021
rect 47578 24012 47584 24024
rect 47636 24012 47642 24064
rect 1104 23962 58880 23984
rect 1104 23910 15398 23962
rect 15450 23910 15462 23962
rect 15514 23910 15526 23962
rect 15578 23910 15590 23962
rect 15642 23910 15654 23962
rect 15706 23910 29846 23962
rect 29898 23910 29910 23962
rect 29962 23910 29974 23962
rect 30026 23910 30038 23962
rect 30090 23910 30102 23962
rect 30154 23910 44294 23962
rect 44346 23910 44358 23962
rect 44410 23910 44422 23962
rect 44474 23910 44486 23962
rect 44538 23910 44550 23962
rect 44602 23910 58880 23962
rect 1104 23888 58880 23910
rect 5810 23848 5816 23860
rect 5460 23820 5816 23848
rect 1581 23783 1639 23789
rect 1581 23749 1593 23783
rect 1627 23780 1639 23783
rect 2958 23780 2964 23792
rect 1627 23752 2964 23780
rect 1627 23749 1639 23752
rect 1581 23743 1639 23749
rect 2958 23740 2964 23752
rect 3016 23780 3022 23792
rect 5460 23789 5488 23820
rect 5810 23808 5816 23820
rect 5868 23808 5874 23860
rect 9030 23808 9036 23860
rect 9088 23848 9094 23860
rect 9306 23848 9312 23860
rect 9088 23820 9312 23848
rect 9088 23808 9094 23820
rect 9306 23808 9312 23820
rect 9364 23808 9370 23860
rect 15194 23848 15200 23860
rect 15155 23820 15200 23848
rect 15194 23808 15200 23820
rect 15252 23808 15258 23860
rect 21177 23851 21235 23857
rect 21177 23817 21189 23851
rect 21223 23848 21235 23851
rect 22462 23848 22468 23860
rect 21223 23820 22468 23848
rect 21223 23817 21235 23820
rect 21177 23811 21235 23817
rect 22462 23808 22468 23820
rect 22520 23848 22526 23860
rect 24781 23851 24839 23857
rect 24781 23848 24793 23851
rect 22520 23820 24793 23848
rect 22520 23808 22526 23820
rect 24781 23817 24793 23820
rect 24827 23817 24839 23851
rect 24781 23811 24839 23817
rect 25130 23808 25136 23860
rect 25188 23848 25194 23860
rect 30377 23851 30435 23857
rect 30377 23848 30389 23851
rect 25188 23820 30389 23848
rect 25188 23808 25194 23820
rect 30377 23817 30389 23820
rect 30423 23817 30435 23851
rect 30377 23811 30435 23817
rect 31113 23851 31171 23857
rect 31113 23817 31125 23851
rect 31159 23848 31171 23851
rect 31202 23848 31208 23860
rect 31159 23820 31208 23848
rect 31159 23817 31171 23820
rect 31113 23811 31171 23817
rect 31202 23808 31208 23820
rect 31260 23808 31266 23860
rect 47578 23848 47584 23860
rect 32324 23820 47584 23848
rect 5445 23783 5503 23789
rect 3016 23752 4016 23780
rect 3016 23740 3022 23752
rect 3988 23724 4016 23752
rect 5445 23749 5457 23783
rect 5491 23749 5503 23783
rect 5445 23743 5503 23749
rect 5661 23783 5719 23789
rect 5661 23749 5673 23783
rect 5707 23780 5719 23783
rect 6086 23780 6092 23792
rect 5707 23752 6092 23780
rect 5707 23749 5719 23752
rect 5661 23743 5719 23749
rect 6086 23740 6092 23752
rect 6144 23740 6150 23792
rect 13170 23780 13176 23792
rect 12742 23752 13176 23780
rect 13170 23740 13176 23752
rect 13228 23740 13234 23792
rect 14642 23740 14648 23792
rect 14700 23780 14706 23792
rect 16945 23783 17003 23789
rect 16945 23780 16957 23783
rect 14700 23752 16957 23780
rect 14700 23740 14706 23752
rect 16945 23749 16957 23752
rect 16991 23749 17003 23783
rect 24578 23780 24584 23792
rect 24539 23752 24584 23780
rect 16945 23743 17003 23749
rect 2038 23712 2044 23724
rect 1999 23684 2044 23712
rect 2038 23672 2044 23684
rect 2096 23672 2102 23724
rect 3050 23712 3056 23724
rect 3011 23684 3056 23712
rect 3050 23672 3056 23684
rect 3108 23672 3114 23724
rect 3326 23712 3332 23724
rect 3287 23684 3332 23712
rect 3326 23672 3332 23684
rect 3384 23672 3390 23724
rect 3970 23712 3976 23724
rect 3931 23684 3976 23712
rect 3970 23672 3976 23684
rect 4028 23672 4034 23724
rect 4798 23712 4804 23724
rect 4759 23684 4804 23712
rect 4798 23672 4804 23684
rect 4856 23672 4862 23724
rect 6549 23715 6607 23721
rect 6549 23681 6561 23715
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 3881 23647 3939 23653
rect 3881 23613 3893 23647
rect 3927 23613 3939 23647
rect 5994 23644 6000 23656
rect 3881 23607 3939 23613
rect 4356 23616 6000 23644
rect 2777 23579 2835 23585
rect 2777 23545 2789 23579
rect 2823 23576 2835 23579
rect 3234 23576 3240 23588
rect 2823 23548 3240 23576
rect 2823 23545 2835 23548
rect 2777 23539 2835 23545
rect 3234 23536 3240 23548
rect 3292 23576 3298 23588
rect 3896 23576 3924 23607
rect 4356 23585 4384 23616
rect 5994 23604 6000 23616
rect 6052 23604 6058 23656
rect 6564 23644 6592 23675
rect 6638 23672 6644 23724
rect 6696 23712 6702 23724
rect 7009 23715 7067 23721
rect 7009 23712 7021 23715
rect 6696 23684 7021 23712
rect 6696 23672 6702 23684
rect 7009 23681 7021 23684
rect 7055 23681 7067 23715
rect 7009 23675 7067 23681
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 8570 23644 8576 23656
rect 6564 23616 8576 23644
rect 8570 23604 8576 23616
rect 8628 23644 8634 23656
rect 9122 23644 9128 23656
rect 8628 23616 9128 23644
rect 8628 23604 8634 23616
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 10980 23644 11008 23675
rect 13446 23672 13452 23724
rect 13504 23712 13510 23724
rect 13906 23712 13912 23724
rect 13504 23684 13549 23712
rect 13867 23684 13912 23712
rect 13504 23672 13510 23684
rect 13906 23672 13912 23684
rect 13964 23672 13970 23724
rect 16761 23715 16819 23721
rect 16761 23681 16773 23715
rect 16807 23681 16819 23715
rect 16960 23712 16988 23743
rect 24578 23740 24584 23752
rect 24636 23740 24642 23792
rect 28813 23783 28871 23789
rect 25884 23752 28120 23780
rect 17957 23715 18015 23721
rect 17957 23712 17969 23715
rect 16960 23684 17969 23712
rect 16761 23675 16819 23681
rect 17957 23681 17969 23684
rect 18003 23712 18015 23715
rect 18322 23712 18328 23724
rect 18003 23684 18328 23712
rect 18003 23681 18015 23684
rect 17957 23675 18015 23681
rect 13078 23644 13084 23656
rect 10980 23616 13084 23644
rect 13078 23604 13084 23616
rect 13136 23604 13142 23656
rect 13173 23647 13231 23653
rect 13173 23613 13185 23647
rect 13219 23644 13231 23647
rect 16114 23644 16120 23656
rect 13219 23616 16120 23644
rect 13219 23613 13231 23616
rect 13173 23607 13231 23613
rect 16114 23604 16120 23616
rect 16172 23604 16178 23656
rect 3292 23548 3924 23576
rect 4341 23579 4399 23585
rect 3292 23536 3298 23548
rect 4341 23545 4353 23579
rect 4387 23545 4399 23579
rect 4341 23539 4399 23545
rect 4893 23579 4951 23585
rect 4893 23545 4905 23579
rect 4939 23576 4951 23579
rect 6362 23576 6368 23588
rect 4939 23548 6368 23576
rect 4939 23545 4951 23548
rect 4893 23539 4951 23545
rect 6362 23536 6368 23548
rect 6420 23536 6426 23588
rect 7834 23536 7840 23588
rect 7892 23576 7898 23588
rect 8297 23579 8355 23585
rect 8297 23576 8309 23579
rect 7892 23548 8309 23576
rect 7892 23536 7898 23548
rect 8297 23545 8309 23548
rect 8343 23545 8355 23579
rect 8297 23539 8355 23545
rect 13446 23536 13452 23588
rect 13504 23576 13510 23588
rect 13722 23576 13728 23588
rect 13504 23548 13728 23576
rect 13504 23536 13510 23548
rect 13722 23536 13728 23548
rect 13780 23536 13786 23588
rect 2222 23508 2228 23520
rect 2183 23480 2228 23508
rect 2222 23468 2228 23480
rect 2280 23468 2286 23520
rect 3145 23511 3203 23517
rect 3145 23477 3157 23511
rect 3191 23508 3203 23511
rect 4154 23508 4160 23520
rect 3191 23480 4160 23508
rect 3191 23477 3203 23480
rect 3145 23471 3203 23477
rect 4154 23468 4160 23480
rect 4212 23468 4218 23520
rect 5626 23508 5632 23520
rect 5587 23480 5632 23508
rect 5626 23468 5632 23480
rect 5684 23468 5690 23520
rect 5810 23508 5816 23520
rect 5771 23480 5816 23508
rect 5810 23468 5816 23480
rect 5868 23468 5874 23520
rect 6457 23511 6515 23517
rect 6457 23477 6469 23511
rect 6503 23508 6515 23511
rect 8018 23508 8024 23520
rect 6503 23480 8024 23508
rect 6503 23477 6515 23480
rect 6457 23471 6515 23477
rect 8018 23468 8024 23480
rect 8076 23468 8082 23520
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 11701 23511 11759 23517
rect 9732 23480 9777 23508
rect 9732 23468 9738 23480
rect 11701 23477 11713 23511
rect 11747 23508 11759 23511
rect 16776 23508 16804 23675
rect 18322 23672 18328 23684
rect 18380 23672 18386 23724
rect 19245 23715 19303 23721
rect 19245 23681 19257 23715
rect 19291 23712 19303 23715
rect 21085 23715 21143 23721
rect 19291 23684 21036 23712
rect 19291 23681 19303 23684
rect 19245 23675 19303 23681
rect 17310 23604 17316 23656
rect 17368 23644 17374 23656
rect 17589 23647 17647 23653
rect 17589 23644 17601 23647
rect 17368 23616 17601 23644
rect 17368 23604 17374 23616
rect 17589 23613 17601 23616
rect 17635 23613 17647 23647
rect 17589 23607 17647 23613
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 19610 23644 19616 23656
rect 18095 23616 19616 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 17604 23576 17632 23607
rect 19610 23604 19616 23616
rect 19668 23604 19674 23656
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23613 19763 23647
rect 19978 23644 19984 23656
rect 19939 23616 19984 23644
rect 19705 23607 19763 23613
rect 19720 23576 19748 23607
rect 19978 23604 19984 23616
rect 20036 23604 20042 23656
rect 21008 23644 21036 23684
rect 21085 23681 21097 23715
rect 21131 23712 21143 23715
rect 21174 23712 21180 23724
rect 21131 23684 21180 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 21174 23672 21180 23684
rect 21232 23672 21238 23724
rect 21269 23715 21327 23721
rect 21269 23681 21281 23715
rect 21315 23712 21327 23715
rect 21910 23712 21916 23724
rect 21315 23684 21916 23712
rect 21315 23681 21327 23684
rect 21269 23675 21327 23681
rect 21910 23672 21916 23684
rect 21968 23672 21974 23724
rect 22002 23672 22008 23724
rect 22060 23712 22066 23724
rect 23293 23715 23351 23721
rect 23293 23712 23305 23715
rect 22060 23684 23305 23712
rect 22060 23672 22066 23684
rect 23293 23681 23305 23684
rect 23339 23681 23351 23715
rect 23293 23675 23351 23681
rect 24394 23672 24400 23724
rect 24452 23712 24458 23724
rect 25884 23721 25912 23752
rect 25869 23715 25927 23721
rect 25869 23712 25881 23715
rect 24452 23684 25881 23712
rect 24452 23672 24458 23684
rect 25869 23681 25881 23684
rect 25915 23681 25927 23715
rect 25869 23675 25927 23681
rect 26418 23672 26424 23724
rect 26476 23712 26482 23724
rect 26970 23712 26976 23724
rect 26476 23684 26976 23712
rect 26476 23672 26482 23684
rect 26970 23672 26976 23684
rect 27028 23712 27034 23724
rect 27065 23715 27123 23721
rect 27065 23712 27077 23715
rect 27028 23684 27077 23712
rect 27028 23672 27034 23684
rect 27065 23681 27077 23684
rect 27111 23681 27123 23715
rect 27982 23712 27988 23724
rect 27943 23684 27988 23712
rect 27065 23675 27123 23681
rect 27982 23672 27988 23684
rect 28040 23672 28046 23724
rect 28092 23712 28120 23752
rect 28813 23749 28825 23783
rect 28859 23780 28871 23783
rect 32324 23780 32352 23820
rect 47578 23808 47584 23820
rect 47636 23808 47642 23860
rect 28859 23752 32352 23780
rect 28859 23749 28871 23752
rect 28813 23743 28871 23749
rect 33870 23740 33876 23792
rect 33928 23780 33934 23792
rect 33965 23783 34023 23789
rect 33965 23780 33977 23783
rect 33928 23752 33977 23780
rect 33928 23740 33934 23752
rect 33965 23749 33977 23752
rect 34011 23749 34023 23783
rect 35986 23780 35992 23792
rect 35190 23752 35992 23780
rect 33965 23743 34023 23749
rect 35986 23740 35992 23752
rect 36044 23740 36050 23792
rect 37550 23780 37556 23792
rect 37511 23752 37556 23780
rect 37550 23740 37556 23752
rect 37608 23740 37614 23792
rect 40678 23740 40684 23792
rect 40736 23780 40742 23792
rect 47765 23783 47823 23789
rect 47765 23780 47777 23783
rect 40736 23752 47777 23780
rect 40736 23740 40742 23752
rect 47765 23749 47777 23752
rect 47811 23749 47823 23783
rect 47765 23743 47823 23749
rect 28092 23684 29500 23712
rect 29472 23656 29500 23684
rect 29546 23672 29552 23724
rect 29604 23712 29610 23724
rect 29604 23684 29649 23712
rect 29604 23672 29610 23684
rect 29822 23672 29828 23724
rect 29880 23712 29886 23724
rect 30469 23715 30527 23721
rect 30469 23712 30481 23715
rect 29880 23684 30481 23712
rect 29880 23672 29886 23684
rect 30469 23681 30481 23684
rect 30515 23681 30527 23715
rect 30469 23675 30527 23681
rect 31205 23715 31263 23721
rect 31205 23681 31217 23715
rect 31251 23712 31263 23715
rect 31846 23712 31852 23724
rect 31251 23684 31852 23712
rect 31251 23681 31263 23684
rect 31205 23675 31263 23681
rect 31846 23672 31852 23684
rect 31904 23672 31910 23724
rect 32125 23715 32183 23721
rect 32125 23681 32137 23715
rect 32171 23712 32183 23715
rect 32674 23712 32680 23724
rect 32171 23684 32680 23712
rect 32171 23681 32183 23684
rect 32125 23675 32183 23681
rect 32674 23672 32680 23684
rect 32732 23672 32738 23724
rect 38654 23672 38660 23724
rect 38712 23672 38718 23724
rect 39114 23672 39120 23724
rect 39172 23712 39178 23724
rect 39761 23715 39819 23721
rect 39761 23712 39773 23715
rect 39172 23684 39773 23712
rect 39172 23672 39178 23684
rect 39761 23681 39773 23684
rect 39807 23681 39819 23715
rect 39761 23675 39819 23681
rect 56594 23672 56600 23724
rect 56652 23712 56658 23724
rect 57885 23715 57943 23721
rect 57885 23712 57897 23715
rect 56652 23684 57897 23712
rect 56652 23672 56658 23684
rect 57885 23681 57897 23684
rect 57931 23681 57943 23715
rect 57885 23675 57943 23681
rect 21450 23644 21456 23656
rect 21008 23616 21456 23644
rect 21450 23604 21456 23616
rect 21508 23644 21514 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21508 23616 21833 23644
rect 21508 23604 21514 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 22097 23647 22155 23653
rect 22097 23613 22109 23647
rect 22143 23613 22155 23647
rect 22097 23607 22155 23613
rect 23569 23647 23627 23653
rect 23569 23613 23581 23647
rect 23615 23644 23627 23647
rect 24486 23644 24492 23656
rect 23615 23616 24492 23644
rect 23615 23613 23627 23616
rect 23569 23607 23627 23613
rect 17604 23548 19748 23576
rect 20254 23536 20260 23588
rect 20312 23576 20318 23588
rect 22112 23576 22140 23607
rect 24486 23604 24492 23616
rect 24544 23604 24550 23656
rect 25498 23604 25504 23656
rect 25556 23644 25562 23656
rect 25593 23647 25651 23653
rect 25593 23644 25605 23647
rect 25556 23616 25605 23644
rect 25556 23604 25562 23616
rect 25593 23613 25605 23616
rect 25639 23613 25651 23647
rect 28074 23644 28080 23656
rect 28035 23616 28080 23644
rect 25593 23607 25651 23613
rect 28074 23604 28080 23616
rect 28132 23604 28138 23656
rect 29270 23644 29276 23656
rect 29231 23616 29276 23644
rect 29270 23604 29276 23616
rect 29328 23604 29334 23656
rect 29454 23644 29460 23656
rect 29415 23616 29460 23644
rect 29454 23604 29460 23616
rect 29512 23604 29518 23656
rect 29638 23644 29644 23656
rect 29599 23616 29644 23644
rect 29638 23604 29644 23616
rect 29696 23604 29702 23656
rect 29733 23647 29791 23653
rect 29733 23613 29745 23647
rect 29779 23613 29791 23647
rect 29733 23607 29791 23613
rect 33689 23647 33747 23653
rect 33689 23613 33701 23647
rect 33735 23613 33747 23647
rect 33689 23607 33747 23613
rect 20312 23548 22140 23576
rect 20312 23536 20318 23548
rect 21836 23520 21864 23548
rect 23382 23536 23388 23588
rect 23440 23576 23446 23588
rect 26602 23576 26608 23588
rect 23440 23548 26608 23576
rect 23440 23536 23446 23548
rect 26602 23536 26608 23548
rect 26660 23536 26666 23588
rect 27249 23579 27307 23585
rect 27249 23545 27261 23579
rect 27295 23576 27307 23579
rect 27522 23576 27528 23588
rect 27295 23548 27528 23576
rect 27295 23545 27307 23548
rect 27249 23539 27307 23545
rect 27522 23536 27528 23548
rect 27580 23576 27586 23588
rect 29748 23576 29776 23607
rect 33704 23576 33732 23607
rect 36538 23604 36544 23656
rect 36596 23644 36602 23656
rect 37277 23647 37335 23653
rect 37277 23644 37289 23647
rect 36596 23616 37289 23644
rect 36596 23604 36602 23616
rect 37277 23613 37289 23616
rect 37323 23613 37335 23647
rect 37277 23607 37335 23613
rect 39025 23647 39083 23653
rect 39025 23613 39037 23647
rect 39071 23644 39083 23647
rect 39669 23647 39727 23653
rect 39669 23644 39681 23647
rect 39071 23616 39681 23644
rect 39071 23613 39083 23616
rect 39025 23607 39083 23613
rect 39669 23613 39681 23616
rect 39715 23644 39727 23647
rect 39850 23644 39856 23656
rect 39715 23616 39856 23644
rect 39715 23613 39727 23616
rect 39669 23607 39727 23613
rect 39850 23604 39856 23616
rect 39908 23604 39914 23656
rect 40589 23647 40647 23653
rect 40589 23613 40601 23647
rect 40635 23644 40647 23647
rect 42702 23644 42708 23656
rect 40635 23616 42708 23644
rect 40635 23613 40647 23616
rect 40589 23607 40647 23613
rect 42702 23604 42708 23616
rect 42760 23604 42766 23656
rect 47486 23604 47492 23656
rect 47544 23644 47550 23656
rect 47581 23647 47639 23653
rect 47581 23644 47593 23647
rect 47544 23616 47593 23644
rect 47544 23604 47550 23616
rect 47581 23613 47593 23616
rect 47627 23613 47639 23647
rect 48590 23644 48596 23656
rect 48551 23616 48596 23644
rect 47581 23607 47639 23613
rect 48590 23604 48596 23616
rect 48648 23604 48654 23656
rect 27580 23548 29776 23576
rect 31726 23548 33732 23576
rect 27580 23536 27586 23548
rect 19150 23508 19156 23520
rect 11747 23480 16804 23508
rect 19111 23480 19156 23508
rect 11747 23477 11759 23480
rect 11701 23471 11759 23477
rect 19150 23468 19156 23480
rect 19208 23468 19214 23520
rect 21818 23468 21824 23520
rect 21876 23468 21882 23520
rect 23566 23468 23572 23520
rect 23624 23508 23630 23520
rect 24118 23508 24124 23520
rect 23624 23480 24124 23508
rect 23624 23468 23630 23480
rect 24118 23468 24124 23480
rect 24176 23468 24182 23520
rect 24670 23468 24676 23520
rect 24728 23508 24734 23520
rect 24765 23511 24823 23517
rect 24765 23508 24777 23511
rect 24728 23480 24777 23508
rect 24728 23468 24734 23480
rect 24765 23477 24777 23480
rect 24811 23477 24823 23511
rect 24765 23471 24823 23477
rect 24949 23511 25007 23517
rect 24949 23477 24961 23511
rect 24995 23508 25007 23511
rect 26050 23508 26056 23520
rect 24995 23480 26056 23508
rect 24995 23477 25007 23480
rect 24949 23471 25007 23477
rect 26050 23468 26056 23480
rect 26108 23468 26114 23520
rect 28718 23468 28724 23520
rect 28776 23508 28782 23520
rect 31726 23508 31754 23548
rect 28776 23480 31754 23508
rect 28776 23468 28782 23480
rect 32122 23468 32128 23520
rect 32180 23508 32186 23520
rect 32217 23511 32275 23517
rect 32217 23508 32229 23511
rect 32180 23480 32229 23508
rect 32180 23468 32186 23480
rect 32217 23477 32229 23480
rect 32263 23477 32275 23511
rect 32217 23471 32275 23477
rect 35437 23511 35495 23517
rect 35437 23477 35449 23511
rect 35483 23508 35495 23511
rect 35894 23508 35900 23520
rect 35483 23480 35900 23508
rect 35483 23477 35495 23480
rect 35437 23471 35495 23477
rect 35894 23468 35900 23480
rect 35952 23468 35958 23520
rect 57882 23468 57888 23520
rect 57940 23508 57946 23520
rect 58069 23511 58127 23517
rect 58069 23508 58081 23511
rect 57940 23480 58081 23508
rect 57940 23468 57946 23480
rect 58069 23477 58081 23480
rect 58115 23477 58127 23511
rect 58069 23471 58127 23477
rect 1104 23418 58880 23440
rect 1104 23366 8174 23418
rect 8226 23366 8238 23418
rect 8290 23366 8302 23418
rect 8354 23366 8366 23418
rect 8418 23366 8430 23418
rect 8482 23366 22622 23418
rect 22674 23366 22686 23418
rect 22738 23366 22750 23418
rect 22802 23366 22814 23418
rect 22866 23366 22878 23418
rect 22930 23366 37070 23418
rect 37122 23366 37134 23418
rect 37186 23366 37198 23418
rect 37250 23366 37262 23418
rect 37314 23366 37326 23418
rect 37378 23366 51518 23418
rect 51570 23366 51582 23418
rect 51634 23366 51646 23418
rect 51698 23366 51710 23418
rect 51762 23366 51774 23418
rect 51826 23366 58880 23418
rect 1104 23344 58880 23366
rect 3970 23264 3976 23316
rect 4028 23304 4034 23316
rect 4028 23276 6684 23304
rect 4028 23264 4034 23276
rect 2685 23239 2743 23245
rect 2685 23205 2697 23239
rect 2731 23236 2743 23239
rect 2866 23236 2872 23248
rect 2731 23208 2872 23236
rect 2731 23205 2743 23208
rect 2685 23199 2743 23205
rect 2866 23196 2872 23208
rect 2924 23196 2930 23248
rect 1581 23171 1639 23177
rect 1581 23137 1593 23171
rect 1627 23168 1639 23171
rect 3145 23171 3203 23177
rect 1627 23140 2268 23168
rect 1627 23137 1639 23140
rect 1581 23131 1639 23137
rect 2240 23112 2268 23140
rect 3145 23137 3157 23171
rect 3191 23168 3203 23171
rect 3234 23168 3240 23180
rect 3191 23140 3240 23168
rect 3191 23137 3203 23140
rect 3145 23131 3203 23137
rect 3234 23128 3240 23140
rect 3292 23128 3298 23180
rect 4157 23171 4215 23177
rect 4157 23137 4169 23171
rect 4203 23168 4215 23171
rect 4522 23168 4528 23180
rect 4203 23140 4528 23168
rect 4203 23137 4215 23140
rect 4157 23131 4215 23137
rect 4522 23128 4528 23140
rect 4580 23128 4586 23180
rect 6546 23168 6552 23180
rect 6507 23140 6552 23168
rect 6546 23128 6552 23140
rect 6604 23128 6610 23180
rect 6656 23168 6684 23276
rect 7558 23264 7564 23316
rect 7616 23304 7622 23316
rect 8297 23307 8355 23313
rect 8297 23304 8309 23307
rect 7616 23276 8309 23304
rect 7616 23264 7622 23276
rect 8297 23273 8309 23276
rect 8343 23273 8355 23307
rect 9858 23304 9864 23316
rect 9819 23276 9864 23304
rect 8297 23267 8355 23273
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 13541 23307 13599 23313
rect 13541 23273 13553 23307
rect 13587 23304 13599 23307
rect 15378 23304 15384 23316
rect 13587 23276 15384 23304
rect 13587 23273 13599 23276
rect 13541 23267 13599 23273
rect 15378 23264 15384 23276
rect 15436 23264 15442 23316
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 18322 23304 18328 23316
rect 18104 23276 18328 23304
rect 18104 23264 18110 23276
rect 18322 23264 18328 23276
rect 18380 23264 18386 23316
rect 18598 23264 18604 23316
rect 18656 23304 18662 23316
rect 18693 23307 18751 23313
rect 18693 23304 18705 23307
rect 18656 23276 18705 23304
rect 18656 23264 18662 23276
rect 18693 23273 18705 23276
rect 18739 23304 18751 23307
rect 19518 23304 19524 23316
rect 18739 23276 19524 23304
rect 18739 23273 18751 23276
rect 18693 23267 18751 23273
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 19797 23307 19855 23313
rect 19797 23273 19809 23307
rect 19843 23304 19855 23307
rect 22186 23304 22192 23316
rect 19843 23276 21036 23304
rect 22099 23276 22192 23304
rect 19843 23273 19855 23276
rect 19797 23267 19855 23273
rect 17034 23236 17040 23248
rect 15764 23208 17040 23236
rect 11146 23168 11152 23180
rect 6656 23140 11152 23168
rect 11146 23128 11152 23140
rect 11204 23128 11210 23180
rect 13630 23168 13636 23180
rect 11348 23140 13636 23168
rect 2038 23100 2044 23112
rect 1999 23072 2044 23100
rect 2038 23060 2044 23072
rect 2096 23060 2102 23112
rect 2222 23060 2228 23112
rect 2280 23100 2286 23112
rect 3053 23103 3111 23109
rect 3053 23100 3065 23103
rect 2280 23072 3065 23100
rect 2280 23060 2286 23072
rect 3053 23069 3065 23072
rect 3099 23069 3111 23103
rect 3878 23100 3884 23112
rect 3839 23072 3884 23100
rect 3053 23063 3111 23069
rect 2225 22967 2283 22973
rect 2225 22933 2237 22967
rect 2271 22964 2283 22967
rect 2774 22964 2780 22976
rect 2271 22936 2780 22964
rect 2271 22933 2283 22936
rect 2225 22927 2283 22933
rect 2774 22924 2780 22936
rect 2832 22924 2838 22976
rect 3068 22964 3096 23063
rect 3878 23060 3884 23072
rect 3936 23060 3942 23112
rect 9125 23103 9183 23109
rect 9125 23069 9137 23103
rect 9171 23100 9183 23103
rect 9674 23100 9680 23112
rect 9171 23072 9680 23100
rect 9171 23069 9183 23072
rect 9125 23063 9183 23069
rect 9674 23060 9680 23072
rect 9732 23100 9738 23112
rect 11054 23100 11060 23112
rect 9732 23072 11060 23100
rect 9732 23060 9738 23072
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 11348 23109 11376 23140
rect 13630 23128 13636 23140
rect 13688 23128 13694 23180
rect 15764 23168 15792 23208
rect 17034 23196 17040 23208
rect 17092 23196 17098 23248
rect 17218 23236 17224 23248
rect 17179 23208 17224 23236
rect 17218 23196 17224 23208
rect 17276 23196 17282 23248
rect 19426 23236 19432 23248
rect 18340 23208 19432 23236
rect 14016 23140 15792 23168
rect 15841 23171 15899 23177
rect 11333 23103 11391 23109
rect 11333 23069 11345 23103
rect 11379 23069 11391 23103
rect 11790 23100 11796 23112
rect 11751 23072 11796 23100
rect 11333 23063 11391 23069
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 13170 23060 13176 23112
rect 13228 23060 13234 23112
rect 4614 22992 4620 23044
rect 4672 22992 4678 23044
rect 6822 23032 6828 23044
rect 5460 23004 5764 23032
rect 6783 23004 6828 23032
rect 5460 22964 5488 23004
rect 3068 22936 5488 22964
rect 5534 22924 5540 22976
rect 5592 22964 5598 22976
rect 5629 22967 5687 22973
rect 5629 22964 5641 22967
rect 5592 22936 5641 22964
rect 5592 22924 5598 22936
rect 5629 22933 5641 22936
rect 5675 22933 5687 22967
rect 5736 22964 5764 23004
rect 6822 22992 6828 23004
rect 6880 22992 6886 23044
rect 7558 22992 7564 23044
rect 7616 22992 7622 23044
rect 12069 23035 12127 23041
rect 8956 23004 10272 23032
rect 8956 22964 8984 23004
rect 5736 22936 8984 22964
rect 9033 22967 9091 22973
rect 5629 22927 5687 22933
rect 9033 22933 9045 22967
rect 9079 22964 9091 22967
rect 10134 22964 10140 22976
rect 9079 22936 10140 22964
rect 9079 22933 9091 22936
rect 9033 22927 9091 22933
rect 10134 22924 10140 22936
rect 10192 22924 10198 22976
rect 10244 22964 10272 23004
rect 12069 23001 12081 23035
rect 12115 23032 12127 23035
rect 12158 23032 12164 23044
rect 12115 23004 12164 23032
rect 12115 23001 12127 23004
rect 12069 22995 12127 23001
rect 12158 22992 12164 23004
rect 12216 22992 12222 23044
rect 14016 22964 14044 23140
rect 15841 23137 15853 23171
rect 15887 23168 15899 23171
rect 15930 23168 15936 23180
rect 15887 23140 15936 23168
rect 15887 23137 15899 23140
rect 15841 23131 15899 23137
rect 15930 23128 15936 23140
rect 15988 23128 15994 23180
rect 18340 23168 18368 23208
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 19536 23236 19564 23264
rect 20901 23239 20959 23245
rect 20901 23236 20913 23239
rect 19536 23208 20913 23236
rect 20901 23205 20913 23208
rect 20947 23205 20959 23239
rect 21008 23236 21036 23276
rect 22186 23264 22192 23276
rect 22244 23304 22250 23316
rect 27430 23304 27436 23316
rect 22244 23276 26740 23304
rect 27391 23276 27436 23304
rect 22244 23264 22250 23276
rect 21008 23208 22094 23236
rect 20901 23199 20959 23205
rect 16500 23140 18368 23168
rect 18417 23171 18475 23177
rect 16500 23109 16528 23140
rect 18417 23137 18429 23171
rect 18463 23168 18475 23171
rect 18874 23168 18880 23180
rect 18463 23140 18880 23168
rect 18463 23137 18475 23140
rect 18417 23131 18475 23137
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 19518 23128 19524 23180
rect 19576 23168 19582 23180
rect 20070 23168 20076 23180
rect 19576 23140 20076 23168
rect 19576 23128 19582 23140
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 20990 23168 20996 23180
rect 20951 23140 20996 23168
rect 20990 23128 20996 23140
rect 21048 23128 21054 23180
rect 22066 23168 22094 23208
rect 22370 23196 22376 23248
rect 22428 23236 22434 23248
rect 22649 23239 22707 23245
rect 22649 23236 22661 23239
rect 22428 23208 22661 23236
rect 22428 23196 22434 23208
rect 22649 23205 22661 23208
rect 22695 23205 22707 23239
rect 22649 23199 22707 23205
rect 23934 23196 23940 23248
rect 23992 23236 23998 23248
rect 24765 23239 24823 23245
rect 24765 23236 24777 23239
rect 23992 23208 24777 23236
rect 23992 23196 23998 23208
rect 24765 23205 24777 23208
rect 24811 23205 24823 23239
rect 26513 23239 26571 23245
rect 24765 23199 24823 23205
rect 24872 23208 26096 23236
rect 23566 23168 23572 23180
rect 22066 23140 23572 23168
rect 23566 23128 23572 23140
rect 23624 23128 23630 23180
rect 23676 23140 24808 23168
rect 16485 23103 16543 23109
rect 16485 23069 16497 23103
rect 16531 23069 16543 23103
rect 16485 23063 16543 23069
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23069 17279 23103
rect 17402 23100 17408 23112
rect 17363 23072 17408 23100
rect 17221 23063 17279 23069
rect 15010 22992 15016 23044
rect 15068 22992 15074 23044
rect 15565 23035 15623 23041
rect 15565 23001 15577 23035
rect 15611 23032 15623 23035
rect 16206 23032 16212 23044
rect 15611 23004 16212 23032
rect 15611 23001 15623 23004
rect 15565 22995 15623 23001
rect 16206 22992 16212 23004
rect 16264 22992 16270 23044
rect 10244 22936 14044 22964
rect 14093 22967 14151 22973
rect 14093 22933 14105 22967
rect 14139 22964 14151 22967
rect 16298 22964 16304 22976
rect 14139 22936 16304 22964
rect 14139 22933 14151 22936
rect 14093 22927 14151 22933
rect 16298 22924 16304 22936
rect 16356 22924 16362 22976
rect 16393 22967 16451 22973
rect 16393 22933 16405 22967
rect 16439 22964 16451 22967
rect 16758 22964 16764 22976
rect 16439 22936 16764 22964
rect 16439 22933 16451 22936
rect 16393 22927 16451 22933
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 17236 22964 17264 23063
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23100 18567 23103
rect 18966 23100 18972 23112
rect 18555 23072 18972 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 19978 23060 19984 23112
rect 20036 23100 20042 23112
rect 20438 23100 20444 23112
rect 20036 23072 20444 23100
rect 20036 23060 20042 23072
rect 20438 23060 20444 23072
rect 20496 23100 20502 23112
rect 20625 23103 20683 23109
rect 20625 23100 20637 23103
rect 20496 23072 20637 23100
rect 20496 23060 20502 23072
rect 20625 23069 20637 23072
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 20772 23103 20830 23109
rect 20772 23069 20784 23103
rect 20818 23100 20830 23103
rect 21174 23100 21180 23112
rect 20818 23072 21180 23100
rect 20818 23069 20830 23072
rect 20772 23063 20830 23069
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 21634 23060 21640 23112
rect 21692 23100 21698 23112
rect 23676 23109 23704 23140
rect 22005 23103 22063 23109
rect 22005 23100 22017 23103
rect 21692 23072 22017 23100
rect 21692 23060 21698 23072
rect 22005 23069 22017 23072
rect 22051 23069 22063 23103
rect 23661 23103 23719 23109
rect 22005 23063 22063 23069
rect 22756 23072 23612 23100
rect 17589 23035 17647 23041
rect 17589 23001 17601 23035
rect 17635 23032 17647 23035
rect 17954 23032 17960 23044
rect 17635 23004 17960 23032
rect 17635 23001 17647 23004
rect 17589 22995 17647 23001
rect 17954 22992 17960 23004
rect 18012 22992 18018 23044
rect 18046 22992 18052 23044
rect 18104 23032 18110 23044
rect 19242 23032 19248 23044
rect 18104 23004 18149 23032
rect 18616 23004 19248 23032
rect 18104 22992 18110 23004
rect 18616 22964 18644 23004
rect 19242 22992 19248 23004
rect 19300 22992 19306 23044
rect 19702 23032 19708 23044
rect 19663 23004 19708 23032
rect 19702 22992 19708 23004
rect 19760 22992 19766 23044
rect 21358 23032 21364 23044
rect 21319 23004 21364 23032
rect 21358 22992 21364 23004
rect 21416 22992 21422 23044
rect 21821 23035 21879 23041
rect 21821 23001 21833 23035
rect 21867 23001 21879 23035
rect 22020 23032 22048 23063
rect 22756 23032 22784 23072
rect 22020 23004 22784 23032
rect 22833 23035 22891 23041
rect 21821 22995 21879 23001
rect 22833 23001 22845 23035
rect 22879 23001 22891 23035
rect 23474 23032 23480 23044
rect 23435 23004 23480 23032
rect 22833 22995 22891 23001
rect 17236 22936 18644 22964
rect 20530 22924 20536 22976
rect 20588 22964 20594 22976
rect 21836 22964 21864 22995
rect 20588 22936 21864 22964
rect 22848 22964 22876 22995
rect 23474 22992 23480 23004
rect 23532 22992 23538 23044
rect 23584 23032 23612 23072
rect 23661 23069 23673 23103
rect 23707 23069 23719 23103
rect 24578 23100 24584 23112
rect 23661 23063 23719 23069
rect 23768 23072 24584 23100
rect 23768 23032 23796 23072
rect 24578 23060 24584 23072
rect 24636 23060 24642 23112
rect 24673 23103 24731 23109
rect 24673 23069 24685 23103
rect 24719 23069 24731 23103
rect 24673 23063 24731 23069
rect 23584 23004 23796 23032
rect 23845 23035 23903 23041
rect 23845 23001 23857 23035
rect 23891 23001 23903 23035
rect 23845 22995 23903 23001
rect 23566 22964 23572 22976
rect 22848 22936 23572 22964
rect 20588 22924 20594 22936
rect 23566 22924 23572 22936
rect 23624 22924 23630 22976
rect 23860 22964 23888 22995
rect 24486 22992 24492 23044
rect 24544 23032 24550 23044
rect 24688 23032 24716 23063
rect 24544 23004 24716 23032
rect 24780 23032 24808 23140
rect 24872 23109 24900 23208
rect 25590 23128 25596 23180
rect 25648 23168 25654 23180
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 25648 23140 25973 23168
rect 25648 23128 25654 23140
rect 25961 23137 25973 23140
rect 26007 23137 26019 23171
rect 26068 23168 26096 23208
rect 26513 23205 26525 23239
rect 26559 23205 26571 23239
rect 26513 23199 26571 23205
rect 26528 23168 26556 23199
rect 26712 23177 26740 23276
rect 27430 23264 27436 23276
rect 27488 23304 27494 23316
rect 27614 23304 27620 23316
rect 27488 23276 27620 23304
rect 27488 23264 27494 23276
rect 27614 23264 27620 23276
rect 27672 23264 27678 23316
rect 33962 23304 33968 23316
rect 33923 23276 33968 23304
rect 33962 23264 33968 23276
rect 34020 23264 34026 23316
rect 35986 23304 35992 23316
rect 35947 23276 35992 23304
rect 35986 23264 35992 23276
rect 36044 23264 36050 23316
rect 38197 23307 38255 23313
rect 38197 23273 38209 23307
rect 38243 23304 38255 23307
rect 38654 23304 38660 23316
rect 38243 23276 38660 23304
rect 38243 23273 38255 23276
rect 38197 23267 38255 23273
rect 38654 23264 38660 23276
rect 38712 23264 38718 23316
rect 28074 23236 28080 23248
rect 28035 23208 28080 23236
rect 28074 23196 28080 23208
rect 28132 23196 28138 23248
rect 26068 23140 26556 23168
rect 26697 23171 26755 23177
rect 25961 23131 26019 23137
rect 26697 23137 26709 23171
rect 26743 23137 26755 23171
rect 28626 23168 28632 23180
rect 26697 23131 26755 23137
rect 26896 23140 28632 23168
rect 26896 23112 26924 23140
rect 28626 23128 28632 23140
rect 28684 23128 28690 23180
rect 31846 23128 31852 23180
rect 31904 23168 31910 23180
rect 36262 23168 36268 23180
rect 31904 23140 36268 23168
rect 31904 23128 31910 23140
rect 24857 23103 24915 23109
rect 24857 23069 24869 23103
rect 24903 23069 24915 23103
rect 24857 23063 24915 23069
rect 24946 23060 24952 23112
rect 25004 23100 25010 23112
rect 25041 23103 25099 23109
rect 25041 23100 25053 23103
rect 25004 23072 25053 23100
rect 25004 23060 25010 23072
rect 25041 23069 25053 23072
rect 25087 23069 25099 23103
rect 25682 23100 25688 23112
rect 25643 23072 25688 23100
rect 25041 23063 25099 23069
rect 25682 23060 25688 23072
rect 25740 23060 25746 23112
rect 25774 23060 25780 23112
rect 25832 23100 25838 23112
rect 26053 23103 26111 23109
rect 25832 23072 25877 23100
rect 25832 23060 25838 23072
rect 26053 23069 26065 23103
rect 26099 23100 26111 23103
rect 26418 23100 26424 23112
rect 26099 23072 26424 23100
rect 26099 23069 26111 23072
rect 26053 23063 26111 23069
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 26602 23060 26608 23112
rect 26660 23100 26666 23112
rect 26878 23100 26884 23112
rect 26660 23072 26753 23100
rect 26839 23072 26884 23100
rect 26660 23060 26666 23072
rect 26878 23060 26884 23072
rect 26936 23060 26942 23112
rect 26970 23060 26976 23112
rect 27028 23100 27034 23112
rect 28166 23100 28172 23112
rect 27028 23072 27073 23100
rect 27172 23072 28172 23100
rect 27028 23060 27034 23072
rect 25501 23035 25559 23041
rect 25501 23032 25513 23035
rect 24780 23004 25513 23032
rect 24544 22992 24550 23004
rect 25501 23001 25513 23004
rect 25547 23001 25559 23035
rect 26620 23032 26648 23060
rect 27172 23032 27200 23072
rect 28166 23060 28172 23072
rect 28224 23060 28230 23112
rect 28994 23060 29000 23112
rect 29052 23100 29058 23112
rect 34072 23109 34100 23140
rect 36262 23128 36268 23140
rect 36320 23168 36326 23180
rect 42518 23168 42524 23180
rect 36320 23140 38148 23168
rect 42479 23140 42524 23168
rect 36320 23128 36326 23140
rect 29549 23103 29607 23109
rect 29549 23100 29561 23103
rect 29052 23072 29561 23100
rect 29052 23060 29058 23072
rect 29549 23069 29561 23072
rect 29595 23069 29607 23103
rect 29549 23063 29607 23069
rect 29825 23103 29883 23109
rect 29825 23069 29837 23103
rect 29871 23100 29883 23103
rect 31113 23103 31171 23109
rect 31113 23100 31125 23103
rect 29871 23072 31125 23100
rect 29871 23069 29883 23072
rect 29825 23063 29883 23069
rect 31113 23069 31125 23072
rect 31159 23069 31171 23103
rect 31113 23063 31171 23069
rect 34057 23103 34115 23109
rect 34057 23069 34069 23103
rect 34103 23069 34115 23103
rect 35434 23100 35440 23112
rect 35395 23072 35440 23100
rect 34057 23063 34115 23069
rect 26620 23004 27200 23032
rect 25501 22995 25559 23001
rect 27982 22992 27988 23044
rect 28040 23032 28046 23044
rect 28077 23035 28135 23041
rect 28077 23032 28089 23035
rect 28040 23004 28089 23032
rect 28040 22992 28046 23004
rect 28077 23001 28089 23004
rect 28123 23001 28135 23035
rect 29840 23032 29868 23063
rect 35434 23060 35440 23072
rect 35492 23060 35498 23112
rect 36081 23103 36139 23109
rect 36081 23100 36093 23103
rect 35866 23072 36093 23100
rect 31386 23032 31392 23044
rect 28077 22995 28135 23001
rect 28184 23004 29868 23032
rect 31347 23004 31392 23032
rect 24397 22967 24455 22973
rect 24397 22964 24409 22967
rect 23860 22936 24409 22964
rect 24397 22933 24409 22936
rect 24443 22964 24455 22967
rect 25130 22964 25136 22976
rect 24443 22936 25136 22964
rect 24443 22933 24455 22936
rect 24397 22927 24455 22933
rect 25130 22924 25136 22936
rect 25188 22924 25194 22976
rect 25774 22924 25780 22976
rect 25832 22964 25838 22976
rect 28184 22964 28212 23004
rect 31386 22992 31392 23004
rect 31444 22992 31450 23044
rect 32122 22992 32128 23044
rect 32180 22992 32186 23044
rect 32674 22992 32680 23044
rect 32732 23032 32738 23044
rect 35866 23032 35894 23072
rect 36081 23069 36093 23072
rect 36127 23100 36139 23103
rect 36354 23100 36360 23112
rect 36127 23072 36360 23100
rect 36127 23069 36139 23072
rect 36081 23063 36139 23069
rect 36354 23060 36360 23072
rect 36412 23060 36418 23112
rect 38120 23109 38148 23140
rect 42518 23128 42524 23140
rect 42576 23128 42582 23180
rect 42702 23128 42708 23180
rect 42760 23168 42766 23180
rect 43165 23171 43223 23177
rect 43165 23168 43177 23171
rect 42760 23140 43177 23168
rect 42760 23128 42766 23140
rect 43165 23137 43177 23140
rect 43211 23137 43223 23171
rect 43165 23131 43223 23137
rect 47578 23128 47584 23180
rect 47636 23168 47642 23180
rect 47949 23171 48007 23177
rect 47949 23168 47961 23171
rect 47636 23140 47961 23168
rect 47636 23128 47642 23140
rect 47949 23137 47961 23140
rect 47995 23137 48007 23171
rect 48590 23168 48596 23180
rect 48551 23140 48596 23168
rect 47949 23131 48007 23137
rect 48590 23128 48596 23140
rect 48648 23128 48654 23180
rect 38105 23103 38163 23109
rect 38105 23069 38117 23103
rect 38151 23100 38163 23103
rect 38378 23100 38384 23112
rect 38151 23072 38384 23100
rect 38151 23069 38163 23072
rect 38105 23063 38163 23069
rect 38378 23060 38384 23072
rect 38436 23060 38442 23112
rect 43346 23060 43352 23112
rect 43404 23100 43410 23112
rect 47762 23100 47768 23112
rect 43404 23072 43449 23100
rect 47723 23072 47768 23100
rect 43404 23060 43410 23072
rect 47762 23060 47768 23072
rect 47820 23060 47826 23112
rect 32732 23004 35894 23032
rect 32732 22992 32738 23004
rect 28534 22964 28540 22976
rect 25832 22936 28212 22964
rect 28495 22936 28540 22964
rect 25832 22924 25838 22936
rect 28534 22924 28540 22936
rect 28592 22924 28598 22976
rect 28810 22964 28816 22976
rect 28771 22936 28816 22964
rect 28810 22924 28816 22936
rect 28868 22924 28874 22976
rect 32858 22964 32864 22976
rect 32819 22936 32864 22964
rect 32858 22924 32864 22936
rect 32916 22924 32922 22976
rect 35066 22924 35072 22976
rect 35124 22964 35130 22976
rect 35345 22967 35403 22973
rect 35345 22964 35357 22967
rect 35124 22936 35357 22964
rect 35124 22924 35130 22936
rect 35345 22933 35357 22936
rect 35391 22933 35403 22967
rect 35345 22927 35403 22933
rect 46201 22967 46259 22973
rect 46201 22933 46213 22967
rect 46247 22964 46259 22967
rect 46566 22964 46572 22976
rect 46247 22936 46572 22964
rect 46247 22933 46259 22936
rect 46201 22927 46259 22933
rect 46566 22924 46572 22936
rect 46624 22964 46630 22976
rect 46661 22967 46719 22973
rect 46661 22964 46673 22967
rect 46624 22936 46673 22964
rect 46624 22924 46630 22936
rect 46661 22933 46673 22936
rect 46707 22933 46719 22967
rect 46661 22927 46719 22933
rect 47305 22967 47363 22973
rect 47305 22933 47317 22967
rect 47351 22964 47363 22967
rect 47394 22964 47400 22976
rect 47351 22936 47400 22964
rect 47351 22933 47363 22936
rect 47305 22927 47363 22933
rect 47394 22924 47400 22936
rect 47452 22924 47458 22976
rect 1104 22874 58880 22896
rect 1104 22822 15398 22874
rect 15450 22822 15462 22874
rect 15514 22822 15526 22874
rect 15578 22822 15590 22874
rect 15642 22822 15654 22874
rect 15706 22822 29846 22874
rect 29898 22822 29910 22874
rect 29962 22822 29974 22874
rect 30026 22822 30038 22874
rect 30090 22822 30102 22874
rect 30154 22822 44294 22874
rect 44346 22822 44358 22874
rect 44410 22822 44422 22874
rect 44474 22822 44486 22874
rect 44538 22822 44550 22874
rect 44602 22822 58880 22874
rect 1104 22800 58880 22822
rect 4525 22763 4583 22769
rect 4525 22729 4537 22763
rect 4571 22760 4583 22763
rect 6638 22760 6644 22772
rect 4571 22732 6644 22760
rect 4571 22729 4583 22732
rect 4525 22723 4583 22729
rect 6638 22720 6644 22732
rect 6696 22720 6702 22772
rect 6730 22720 6736 22772
rect 6788 22760 6794 22772
rect 6914 22760 6920 22772
rect 6788 22732 6920 22760
rect 6788 22720 6794 22732
rect 6914 22720 6920 22732
rect 6972 22760 6978 22772
rect 7742 22760 7748 22772
rect 6972 22732 7748 22760
rect 6972 22720 6978 22732
rect 7742 22720 7748 22732
rect 7800 22720 7806 22772
rect 8018 22720 8024 22772
rect 8076 22760 8082 22772
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 8076 22732 9260 22760
rect 8076 22720 8082 22732
rect 3050 22692 3056 22704
rect 2148 22664 3056 22692
rect 2148 22633 2176 22664
rect 3050 22652 3056 22664
rect 3108 22652 3114 22704
rect 7006 22692 7012 22704
rect 5828 22664 7012 22692
rect 2133 22627 2191 22633
rect 2133 22593 2145 22627
rect 2179 22593 2191 22627
rect 2133 22587 2191 22593
rect 2685 22627 2743 22633
rect 2685 22593 2697 22627
rect 2731 22624 2743 22627
rect 4341 22627 4399 22633
rect 2731 22596 4292 22624
rect 2731 22593 2743 22596
rect 2685 22587 2743 22593
rect 4264 22556 4292 22596
rect 4341 22593 4353 22627
rect 4387 22624 4399 22627
rect 4706 22624 4712 22636
rect 4387 22596 4712 22624
rect 4387 22593 4399 22596
rect 4341 22587 4399 22593
rect 4706 22584 4712 22596
rect 4764 22624 4770 22636
rect 5828 22633 5856 22664
rect 7006 22652 7012 22664
rect 7064 22652 7070 22704
rect 7650 22652 7656 22704
rect 7708 22652 7714 22704
rect 5169 22627 5227 22633
rect 5169 22624 5181 22627
rect 4764 22596 5181 22624
rect 4764 22584 4770 22596
rect 5169 22593 5181 22596
rect 5215 22593 5227 22627
rect 5169 22587 5227 22593
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22593 5871 22627
rect 5813 22587 5871 22593
rect 6362 22584 6368 22636
rect 6420 22624 6426 22636
rect 9232 22633 9260 22732
rect 9876 22732 13093 22760
rect 9766 22652 9772 22704
rect 9824 22692 9830 22704
rect 9876 22692 9904 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 13081 22723 13139 22729
rect 13262 22720 13268 22772
rect 13320 22760 13326 22772
rect 13722 22760 13728 22772
rect 13320 22732 13728 22760
rect 13320 22720 13326 22732
rect 13722 22720 13728 22732
rect 13780 22720 13786 22772
rect 14918 22720 14924 22772
rect 14976 22760 14982 22772
rect 14976 22732 15148 22760
rect 14976 22720 14982 22732
rect 9824 22664 9982 22692
rect 9824 22652 9830 22664
rect 11054 22652 11060 22704
rect 11112 22692 11118 22704
rect 14090 22692 14096 22704
rect 11112 22664 12572 22692
rect 11112 22652 11118 22664
rect 12544 22636 12572 22664
rect 13740 22664 14096 22692
rect 6733 22628 6791 22633
rect 6656 22627 6791 22628
rect 6656 22624 6745 22627
rect 6420 22600 6745 22624
rect 6420 22596 6684 22600
rect 6420 22584 6426 22596
rect 6733 22593 6745 22600
rect 6779 22593 6791 22627
rect 6733 22587 6791 22593
rect 9217 22627 9275 22633
rect 9217 22593 9229 22627
rect 9263 22593 9275 22627
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 9217 22587 9275 22593
rect 10980 22596 11529 22624
rect 6638 22556 6644 22568
rect 4264 22528 6644 22556
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 7009 22559 7067 22565
rect 7009 22525 7021 22559
rect 7055 22556 7067 22559
rect 7098 22556 7104 22568
rect 7055 22528 7104 22556
rect 7055 22525 7067 22528
rect 7009 22519 7067 22525
rect 7098 22516 7104 22528
rect 7156 22516 7162 22568
rect 7742 22516 7748 22568
rect 7800 22556 7806 22568
rect 10980 22565 11008 22596
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 11517 22587 11575 22593
rect 12526 22584 12532 22636
rect 12584 22622 12590 22636
rect 13170 22624 13176 22636
rect 12584 22594 12627 22622
rect 13131 22596 13176 22624
rect 12584 22584 12590 22594
rect 13170 22584 13176 22596
rect 13228 22584 13234 22636
rect 13740 22633 13768 22664
rect 14090 22652 14096 22664
rect 14148 22652 14154 22704
rect 13725 22627 13783 22633
rect 13725 22593 13737 22627
rect 13771 22593 13783 22627
rect 15120 22610 15148 22732
rect 17034 22720 17040 22772
rect 17092 22760 17098 22772
rect 17310 22760 17316 22772
rect 17092 22732 17316 22760
rect 17092 22720 17098 22732
rect 17310 22720 17316 22732
rect 17368 22760 17374 22772
rect 17405 22763 17463 22769
rect 17405 22760 17417 22763
rect 17368 22732 17417 22760
rect 17368 22720 17374 22732
rect 17405 22729 17417 22732
rect 17451 22729 17463 22763
rect 17405 22723 17463 22729
rect 20809 22763 20867 22769
rect 20809 22729 20821 22763
rect 20855 22760 20867 22763
rect 20898 22760 20904 22772
rect 20855 22732 20904 22760
rect 20855 22729 20867 22732
rect 20809 22723 20867 22729
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 21266 22720 21272 22772
rect 21324 22760 21330 22772
rect 21324 22732 24164 22760
rect 21324 22720 21330 22732
rect 23474 22692 23480 22704
rect 19812 22664 23480 22692
rect 13725 22587 13783 22593
rect 16022 22584 16028 22636
rect 16080 22624 16086 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 16080 22596 16129 22624
rect 16080 22584 16086 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 16117 22587 16175 22593
rect 16298 22584 16304 22636
rect 16356 22624 16362 22636
rect 16669 22627 16727 22633
rect 16669 22624 16681 22627
rect 16356 22596 16681 22624
rect 16356 22584 16362 22596
rect 16669 22593 16681 22596
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 17402 22584 17408 22636
rect 17460 22624 17466 22636
rect 17770 22624 17776 22636
rect 17460 22596 17776 22624
rect 17460 22584 17466 22596
rect 17770 22584 17776 22596
rect 17828 22624 17834 22636
rect 19812 22633 19840 22664
rect 23474 22652 23480 22664
rect 23532 22652 23538 22704
rect 24136 22636 24164 22732
rect 24210 22720 24216 22772
rect 24268 22760 24274 22772
rect 24578 22760 24584 22772
rect 24268 22732 24584 22760
rect 24268 22720 24274 22732
rect 24578 22720 24584 22732
rect 24636 22720 24642 22772
rect 24670 22720 24676 22772
rect 24728 22760 24734 22772
rect 25314 22760 25320 22772
rect 24728 22732 24808 22760
rect 25275 22732 25320 22760
rect 24728 22720 24734 22732
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 17828 22596 18889 22624
rect 17828 22584 17834 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 19797 22627 19855 22633
rect 19797 22593 19809 22627
rect 19843 22593 19855 22627
rect 19797 22587 19855 22593
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 21177 22627 21235 22633
rect 21177 22624 21189 22627
rect 20772 22596 21189 22624
rect 20772 22584 20778 22596
rect 21177 22593 21189 22596
rect 21223 22593 21235 22627
rect 22278 22624 22284 22636
rect 21177 22587 21235 22593
rect 21560 22596 22284 22624
rect 8757 22559 8815 22565
rect 8757 22556 8769 22559
rect 7800 22528 8769 22556
rect 7800 22516 7806 22528
rect 8757 22525 8769 22528
rect 8803 22525 8815 22559
rect 9493 22559 9551 22565
rect 9493 22556 9505 22559
rect 8757 22519 8815 22525
rect 8864 22528 9505 22556
rect 2958 22448 2964 22500
rect 3016 22488 3022 22500
rect 3145 22491 3203 22497
rect 3145 22488 3157 22491
rect 3016 22460 3157 22488
rect 3016 22448 3022 22460
rect 3145 22457 3157 22460
rect 3191 22457 3203 22491
rect 3145 22451 3203 22457
rect 4982 22420 4988 22432
rect 4943 22392 4988 22420
rect 4982 22380 4988 22392
rect 5040 22380 5046 22432
rect 5721 22423 5779 22429
rect 5721 22389 5733 22423
rect 5767 22420 5779 22423
rect 5810 22420 5816 22432
rect 5767 22392 5816 22420
rect 5767 22389 5779 22392
rect 5721 22383 5779 22389
rect 5810 22380 5816 22392
rect 5868 22380 5874 22432
rect 5994 22380 6000 22432
rect 6052 22420 6058 22432
rect 8864 22420 8892 22528
rect 9493 22525 9505 22528
rect 9539 22525 9551 22559
rect 9493 22519 9551 22525
rect 10965 22559 11023 22565
rect 10965 22525 10977 22559
rect 11011 22525 11023 22559
rect 10965 22519 11023 22525
rect 14001 22559 14059 22565
rect 14001 22525 14013 22559
rect 14047 22556 14059 22559
rect 15286 22556 15292 22568
rect 14047 22528 15292 22556
rect 14047 22525 14059 22528
rect 14001 22519 14059 22525
rect 15286 22516 15292 22528
rect 15344 22516 15350 22568
rect 16574 22516 16580 22568
rect 16632 22556 16638 22568
rect 21085 22559 21143 22565
rect 16632 22528 18552 22556
rect 16632 22516 16638 22528
rect 11146 22448 11152 22500
rect 11204 22488 11210 22500
rect 11701 22491 11759 22497
rect 11701 22488 11713 22491
rect 11204 22460 11713 22488
rect 11204 22448 11210 22460
rect 11701 22457 11713 22460
rect 11747 22488 11759 22491
rect 15473 22491 15531 22497
rect 11747 22460 13492 22488
rect 11747 22457 11759 22460
rect 11701 22451 11759 22457
rect 6052 22392 8892 22420
rect 6052 22380 6058 22392
rect 12434 22380 12440 22432
rect 12492 22420 12498 22432
rect 13464 22420 13492 22460
rect 15473 22457 15485 22491
rect 15519 22488 15531 22491
rect 17126 22488 17132 22500
rect 15519 22460 17132 22488
rect 15519 22457 15531 22460
rect 15473 22451 15531 22457
rect 17126 22448 17132 22460
rect 17184 22448 17190 22500
rect 18414 22488 18420 22500
rect 18375 22460 18420 22488
rect 18414 22448 18420 22460
rect 18472 22448 18478 22500
rect 18524 22488 18552 22528
rect 21085 22525 21097 22559
rect 21131 22556 21143 22559
rect 21560 22556 21588 22596
rect 22278 22584 22284 22596
rect 22336 22584 22342 22636
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 23293 22627 23351 22633
rect 23293 22593 23305 22627
rect 23339 22624 23351 22627
rect 23658 22624 23664 22636
rect 23339 22596 23664 22624
rect 23339 22593 23351 22596
rect 23293 22587 23351 22593
rect 21818 22556 21824 22568
rect 21131 22528 21588 22556
rect 21779 22528 21824 22556
rect 21131 22525 21143 22528
rect 21085 22519 21143 22525
rect 21818 22516 21824 22528
rect 21876 22516 21882 22568
rect 22097 22559 22155 22565
rect 22097 22525 22109 22559
rect 22143 22556 22155 22559
rect 23124 22556 23152 22587
rect 23658 22584 23664 22596
rect 23716 22584 23722 22636
rect 23842 22624 23848 22636
rect 23803 22596 23848 22624
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 24118 22624 24124 22636
rect 24031 22596 24124 22624
rect 24118 22584 24124 22596
rect 24176 22624 24182 22636
rect 24670 22624 24676 22636
rect 24176 22596 24676 22624
rect 24176 22584 24182 22596
rect 24670 22584 24676 22596
rect 24728 22584 24734 22636
rect 24780 22633 24808 22732
rect 25314 22720 25320 22732
rect 25372 22720 25378 22772
rect 25682 22720 25688 22772
rect 25740 22760 25746 22772
rect 26145 22763 26203 22769
rect 26145 22760 26157 22763
rect 25740 22732 26157 22760
rect 25740 22720 25746 22732
rect 26145 22729 26157 22732
rect 26191 22729 26203 22763
rect 26145 22723 26203 22729
rect 31386 22720 31392 22772
rect 31444 22760 31450 22772
rect 32953 22763 33011 22769
rect 32953 22760 32965 22763
rect 31444 22732 32965 22760
rect 31444 22720 31450 22732
rect 32953 22729 32965 22732
rect 32999 22729 33011 22763
rect 32953 22723 33011 22729
rect 44468 22732 47072 22760
rect 25777 22695 25835 22701
rect 25777 22692 25789 22695
rect 25056 22664 25789 22692
rect 24765 22627 24823 22633
rect 24765 22593 24777 22627
rect 24811 22624 24823 22627
rect 24946 22624 24952 22636
rect 24811 22596 24952 22624
rect 24811 22593 24823 22596
rect 24765 22587 24823 22593
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 25056 22633 25084 22664
rect 25777 22661 25789 22664
rect 25823 22661 25835 22695
rect 27982 22692 27988 22704
rect 25777 22655 25835 22661
rect 27264 22664 27988 22692
rect 25041 22627 25099 22633
rect 25041 22593 25053 22627
rect 25087 22593 25099 22627
rect 25041 22587 25099 22593
rect 25130 22584 25136 22636
rect 25188 22624 25194 22636
rect 25188 22596 25233 22624
rect 25188 22584 25194 22596
rect 25498 22584 25504 22636
rect 25556 22624 25562 22636
rect 25961 22627 26019 22633
rect 25961 22624 25973 22627
rect 25556 22596 25973 22624
rect 25556 22584 25562 22596
rect 25961 22593 25973 22596
rect 26007 22593 26019 22627
rect 25961 22587 26019 22593
rect 26234 22584 26240 22636
rect 26292 22624 26298 22636
rect 26292 22596 26337 22624
rect 26292 22584 26298 22596
rect 26418 22584 26424 22636
rect 26476 22624 26482 22636
rect 27264 22633 27292 22664
rect 27982 22652 27988 22664
rect 28040 22652 28046 22704
rect 32217 22695 32275 22701
rect 32217 22692 32229 22695
rect 31326 22664 32229 22692
rect 32217 22661 32229 22664
rect 32263 22661 32275 22695
rect 32217 22655 32275 22661
rect 35066 22652 35072 22704
rect 35124 22652 35130 22704
rect 35529 22695 35587 22701
rect 35529 22661 35541 22695
rect 35575 22692 35587 22695
rect 36357 22695 36415 22701
rect 36357 22692 36369 22695
rect 35575 22664 36369 22692
rect 35575 22661 35587 22664
rect 35529 22655 35587 22661
rect 36357 22661 36369 22664
rect 36403 22661 36415 22695
rect 36357 22655 36415 22661
rect 40681 22695 40739 22701
rect 40681 22661 40693 22695
rect 40727 22692 40739 22695
rect 40770 22692 40776 22704
rect 40727 22664 40776 22692
rect 40727 22661 40739 22664
rect 40681 22655 40739 22661
rect 40770 22652 40776 22664
rect 40828 22652 40834 22704
rect 27249 22627 27307 22633
rect 27249 22624 27261 22627
rect 26476 22596 27261 22624
rect 26476 22584 26482 22596
rect 27249 22593 27261 22596
rect 27295 22593 27307 22627
rect 27249 22587 27307 22593
rect 27433 22627 27491 22633
rect 27433 22593 27445 22627
rect 27479 22593 27491 22627
rect 27433 22587 27491 22593
rect 23934 22556 23940 22568
rect 22143 22528 23152 22556
rect 23895 22528 23940 22556
rect 22143 22525 22155 22528
rect 22097 22519 22155 22525
rect 21266 22488 21272 22500
rect 18524 22460 21272 22488
rect 21266 22448 21272 22460
rect 21324 22448 21330 22500
rect 23124 22488 23152 22528
rect 23934 22516 23940 22528
rect 23992 22516 23998 22568
rect 24857 22559 24915 22565
rect 24857 22525 24869 22559
rect 24903 22556 24915 22559
rect 25590 22556 25596 22568
rect 24903 22528 25596 22556
rect 24903 22525 24915 22528
rect 24857 22519 24915 22525
rect 24210 22488 24216 22500
rect 23124 22460 24216 22488
rect 24210 22448 24216 22460
rect 24268 22448 24274 22500
rect 24305 22491 24363 22497
rect 24305 22457 24317 22491
rect 24351 22488 24363 22491
rect 24872 22488 24900 22519
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 27157 22559 27215 22565
rect 27157 22525 27169 22559
rect 27203 22556 27215 22559
rect 27338 22556 27344 22568
rect 27203 22528 27344 22556
rect 27203 22525 27215 22528
rect 27157 22519 27215 22525
rect 27338 22516 27344 22528
rect 27396 22516 27402 22568
rect 27448 22556 27476 22587
rect 28626 22584 28632 22636
rect 28684 22624 28690 22636
rect 29825 22627 29883 22633
rect 29825 22624 29837 22627
rect 28684 22596 29837 22624
rect 28684 22584 28690 22596
rect 29825 22593 29837 22596
rect 29871 22593 29883 22627
rect 29825 22587 29883 22593
rect 31846 22584 31852 22636
rect 31904 22624 31910 22636
rect 32309 22627 32367 22633
rect 32309 22624 32321 22627
rect 31904 22596 32321 22624
rect 31904 22584 31910 22596
rect 32309 22593 32321 22596
rect 32355 22624 32367 22627
rect 32674 22624 32680 22636
rect 32355 22596 32680 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 32674 22584 32680 22596
rect 32732 22584 32738 22636
rect 33045 22627 33103 22633
rect 33045 22593 33057 22627
rect 33091 22624 33103 22627
rect 33502 22624 33508 22636
rect 33091 22596 33508 22624
rect 33091 22593 33103 22596
rect 33045 22587 33103 22593
rect 33502 22584 33508 22596
rect 33560 22584 33566 22636
rect 35894 22584 35900 22636
rect 35952 22624 35958 22636
rect 36265 22627 36323 22633
rect 36265 22624 36277 22627
rect 35952 22596 36277 22624
rect 35952 22584 35958 22596
rect 36265 22593 36277 22596
rect 36311 22593 36323 22627
rect 37734 22624 37740 22636
rect 37695 22596 37740 22624
rect 36265 22587 36323 22593
rect 37734 22584 37740 22596
rect 37792 22584 37798 22636
rect 38378 22624 38384 22636
rect 38339 22596 38384 22624
rect 38378 22584 38384 22596
rect 38436 22584 38442 22636
rect 39301 22627 39359 22633
rect 39301 22593 39313 22627
rect 39347 22624 39359 22627
rect 39758 22624 39764 22636
rect 39347 22596 39764 22624
rect 39347 22593 39359 22596
rect 39301 22587 39359 22593
rect 39758 22584 39764 22596
rect 39816 22584 39822 22636
rect 40954 22624 40960 22636
rect 40915 22596 40960 22624
rect 40954 22584 40960 22596
rect 41012 22584 41018 22636
rect 41601 22627 41659 22633
rect 41601 22593 41613 22627
rect 41647 22624 41659 22627
rect 42518 22624 42524 22636
rect 41647 22596 42524 22624
rect 41647 22593 41659 22596
rect 41601 22587 41659 22593
rect 42518 22584 42524 22596
rect 42576 22584 42582 22636
rect 43346 22584 43352 22636
rect 43404 22624 43410 22636
rect 44468 22633 44496 22732
rect 45646 22652 45652 22704
rect 45704 22692 45710 22704
rect 45704 22664 46046 22692
rect 45704 22652 45710 22664
rect 44453 22627 44511 22633
rect 44453 22624 44465 22627
rect 43404 22596 44465 22624
rect 43404 22584 43410 22596
rect 44453 22593 44465 22596
rect 44499 22593 44511 22627
rect 44453 22587 44511 22593
rect 28077 22559 28135 22565
rect 28077 22556 28089 22559
rect 27448 22528 28089 22556
rect 24351 22460 24900 22488
rect 24351 22457 24363 22460
rect 24305 22451 24363 22457
rect 24946 22448 24952 22500
rect 25004 22488 25010 22500
rect 25774 22488 25780 22500
rect 25004 22460 25780 22488
rect 25004 22448 25010 22460
rect 25774 22448 25780 22460
rect 25832 22488 25838 22500
rect 26234 22488 26240 22500
rect 25832 22460 26240 22488
rect 25832 22448 25838 22460
rect 26234 22448 26240 22460
rect 26292 22448 26298 22500
rect 14458 22420 14464 22432
rect 12492 22392 12537 22420
rect 13464 22392 14464 22420
rect 12492 22380 12498 22392
rect 14458 22380 14464 22392
rect 14516 22380 14522 22432
rect 16022 22420 16028 22432
rect 15983 22392 16028 22420
rect 16022 22380 16028 22392
rect 16080 22380 16086 22432
rect 16574 22380 16580 22432
rect 16632 22420 16638 22432
rect 16853 22423 16911 22429
rect 16853 22420 16865 22423
rect 16632 22392 16865 22420
rect 16632 22380 16638 22392
rect 16853 22389 16865 22392
rect 16899 22389 16911 22423
rect 16853 22383 16911 22389
rect 18506 22380 18512 22432
rect 18564 22420 18570 22432
rect 20622 22420 20628 22432
rect 18564 22392 20628 22420
rect 18564 22380 18570 22392
rect 20622 22380 20628 22392
rect 20680 22380 20686 22432
rect 21174 22420 21180 22432
rect 21087 22392 21180 22420
rect 21174 22380 21180 22392
rect 21232 22420 21238 22432
rect 23198 22420 23204 22432
rect 21232 22392 23204 22420
rect 21232 22380 21238 22392
rect 23198 22380 23204 22392
rect 23256 22380 23262 22432
rect 23750 22380 23756 22432
rect 23808 22420 23814 22432
rect 23845 22423 23903 22429
rect 23845 22420 23857 22423
rect 23808 22392 23857 22420
rect 23808 22380 23814 22392
rect 23845 22389 23857 22392
rect 23891 22389 23903 22423
rect 23845 22383 23903 22389
rect 24026 22380 24032 22432
rect 24084 22420 24090 22432
rect 27448 22420 27476 22528
rect 28077 22525 28089 22528
rect 28123 22525 28135 22559
rect 28077 22519 28135 22525
rect 28353 22559 28411 22565
rect 28353 22525 28365 22559
rect 28399 22556 28411 22559
rect 30098 22556 30104 22568
rect 28399 22528 29132 22556
rect 30059 22528 30104 22556
rect 28399 22525 28411 22528
rect 28353 22519 28411 22525
rect 29104 22432 29132 22528
rect 30098 22516 30104 22528
rect 30156 22516 30162 22568
rect 35805 22559 35863 22565
rect 35805 22556 35817 22559
rect 31726 22528 35817 22556
rect 31726 22488 31754 22528
rect 35805 22525 35817 22528
rect 35851 22556 35863 22559
rect 36538 22556 36544 22568
rect 35851 22528 36544 22556
rect 35851 22525 35863 22528
rect 35805 22519 35863 22525
rect 36538 22516 36544 22528
rect 36596 22516 36602 22568
rect 41874 22516 41880 22568
rect 41932 22556 41938 22568
rect 44545 22559 44603 22565
rect 41932 22528 41977 22556
rect 41932 22516 41938 22528
rect 44545 22525 44557 22559
rect 44591 22556 44603 22559
rect 45278 22556 45284 22568
rect 44591 22528 44772 22556
rect 45239 22528 45284 22556
rect 44591 22525 44603 22528
rect 44545 22519 44603 22525
rect 31128 22460 31754 22488
rect 24084 22392 27476 22420
rect 27617 22423 27675 22429
rect 24084 22380 24090 22392
rect 27617 22389 27629 22423
rect 27663 22420 27675 22423
rect 27798 22420 27804 22432
rect 27663 22392 27804 22420
rect 27663 22389 27675 22392
rect 27617 22383 27675 22389
rect 27798 22380 27804 22392
rect 27856 22380 27862 22432
rect 29086 22380 29092 22432
rect 29144 22420 29150 22432
rect 29638 22420 29644 22432
rect 29144 22392 29644 22420
rect 29144 22380 29150 22392
rect 29638 22380 29644 22392
rect 29696 22420 29702 22432
rect 31128 22420 31156 22460
rect 31570 22420 31576 22432
rect 29696 22392 31156 22420
rect 31531 22392 31576 22420
rect 29696 22380 29702 22392
rect 31570 22380 31576 22392
rect 31628 22380 31634 22432
rect 34054 22420 34060 22432
rect 34015 22392 34060 22420
rect 34054 22380 34060 22392
rect 34112 22380 34118 22432
rect 37734 22380 37740 22432
rect 37792 22420 37798 22432
rect 37829 22423 37887 22429
rect 37829 22420 37841 22423
rect 37792 22392 37841 22420
rect 37792 22380 37798 22392
rect 37829 22389 37841 22392
rect 37875 22389 37887 22423
rect 37829 22383 37887 22389
rect 38473 22423 38531 22429
rect 38473 22389 38485 22423
rect 38519 22420 38531 22423
rect 38746 22420 38752 22432
rect 38519 22392 38752 22420
rect 38519 22389 38531 22392
rect 38473 22383 38531 22389
rect 38746 22380 38752 22392
rect 38804 22380 38810 22432
rect 39206 22420 39212 22432
rect 39167 22392 39212 22420
rect 39206 22380 39212 22392
rect 39264 22380 39270 22432
rect 42518 22420 42524 22432
rect 42479 22392 42524 22420
rect 42518 22380 42524 22392
rect 42576 22380 42582 22432
rect 44744 22420 44772 22528
rect 45278 22516 45284 22528
rect 45336 22516 45342 22568
rect 45557 22559 45615 22565
rect 45557 22556 45569 22559
rect 45388 22528 45569 22556
rect 44821 22491 44879 22497
rect 44821 22457 44833 22491
rect 44867 22488 44879 22491
rect 45388 22488 45416 22528
rect 45557 22525 45569 22528
rect 45603 22525 45615 22559
rect 45557 22519 45615 22525
rect 44867 22460 45416 22488
rect 44867 22457 44879 22460
rect 44821 22451 44879 22457
rect 46566 22448 46572 22500
rect 46624 22488 46630 22500
rect 47044 22497 47072 22732
rect 48314 22692 48320 22704
rect 48275 22664 48320 22692
rect 48314 22652 48320 22664
rect 48372 22652 48378 22704
rect 50525 22627 50583 22633
rect 50525 22624 50537 22627
rect 49528 22596 50537 22624
rect 47670 22516 47676 22568
rect 47728 22556 47734 22568
rect 48133 22559 48191 22565
rect 48133 22556 48145 22559
rect 47728 22528 48145 22556
rect 47728 22516 47734 22528
rect 48133 22525 48145 22528
rect 48179 22525 48191 22559
rect 48590 22556 48596 22568
rect 48503 22528 48596 22556
rect 48133 22519 48191 22525
rect 48590 22516 48596 22528
rect 48648 22516 48654 22568
rect 49142 22516 49148 22568
rect 49200 22556 49206 22568
rect 49528 22556 49556 22596
rect 50525 22593 50537 22596
rect 50571 22593 50583 22627
rect 50525 22587 50583 22593
rect 51813 22627 51871 22633
rect 51813 22593 51825 22627
rect 51859 22624 51871 22627
rect 51902 22624 51908 22636
rect 51859 22596 51908 22624
rect 51859 22593 51871 22596
rect 51813 22587 51871 22593
rect 51902 22584 51908 22596
rect 51960 22584 51966 22636
rect 49200 22528 49556 22556
rect 49200 22516 49206 22528
rect 47029 22491 47087 22497
rect 46624 22460 46980 22488
rect 46624 22448 46630 22460
rect 46842 22420 46848 22432
rect 44744 22392 46848 22420
rect 46842 22380 46848 22392
rect 46900 22380 46906 22432
rect 46952 22420 46980 22460
rect 47029 22457 47041 22491
rect 47075 22488 47087 22491
rect 48038 22488 48044 22500
rect 47075 22460 48044 22488
rect 47075 22457 47087 22460
rect 47029 22451 47087 22457
rect 48038 22448 48044 22460
rect 48096 22448 48102 22500
rect 47581 22423 47639 22429
rect 47581 22420 47593 22423
rect 46952 22392 47593 22420
rect 47581 22389 47593 22392
rect 47627 22420 47639 22423
rect 48608 22420 48636 22516
rect 50709 22491 50767 22497
rect 50709 22457 50721 22491
rect 50755 22488 50767 22491
rect 52270 22488 52276 22500
rect 50755 22460 52276 22488
rect 50755 22457 50767 22460
rect 50709 22451 50767 22457
rect 52270 22448 52276 22460
rect 52328 22448 52334 22500
rect 51994 22420 52000 22432
rect 47627 22392 48636 22420
rect 51955 22392 52000 22420
rect 47627 22389 47639 22392
rect 47581 22383 47639 22389
rect 51994 22380 52000 22392
rect 52052 22380 52058 22432
rect 1104 22330 58880 22352
rect 1104 22278 8174 22330
rect 8226 22278 8238 22330
rect 8290 22278 8302 22330
rect 8354 22278 8366 22330
rect 8418 22278 8430 22330
rect 8482 22278 22622 22330
rect 22674 22278 22686 22330
rect 22738 22278 22750 22330
rect 22802 22278 22814 22330
rect 22866 22278 22878 22330
rect 22930 22278 37070 22330
rect 37122 22278 37134 22330
rect 37186 22278 37198 22330
rect 37250 22278 37262 22330
rect 37314 22278 37326 22330
rect 37378 22278 51518 22330
rect 51570 22278 51582 22330
rect 51634 22278 51646 22330
rect 51698 22278 51710 22330
rect 51762 22278 51774 22330
rect 51826 22278 58880 22330
rect 1104 22256 58880 22278
rect 4706 22216 4712 22228
rect 4667 22188 4712 22216
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 6886 22188 9444 22216
rect 2317 22151 2375 22157
rect 2317 22117 2329 22151
rect 2363 22148 2375 22151
rect 6886 22148 6914 22188
rect 2363 22120 6914 22148
rect 2363 22117 2375 22120
rect 2317 22111 2375 22117
rect 2041 22083 2099 22089
rect 2041 22049 2053 22083
rect 2087 22080 2099 22083
rect 2222 22080 2228 22092
rect 2087 22052 2228 22080
rect 2087 22049 2099 22052
rect 2041 22043 2099 22049
rect 2222 22040 2228 22052
rect 2280 22040 2286 22092
rect 3881 22083 3939 22089
rect 3881 22049 3893 22083
rect 3927 22080 3939 22083
rect 4614 22080 4620 22092
rect 3927 22052 4620 22080
rect 3927 22049 3939 22052
rect 3881 22043 3939 22049
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 7374 22040 7380 22092
rect 7432 22080 7438 22092
rect 9416 22089 9444 22188
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 13093 22219 13151 22225
rect 13093 22216 13105 22219
rect 11388 22188 13105 22216
rect 11388 22176 11394 22188
rect 13093 22185 13105 22188
rect 13139 22185 13151 22219
rect 13093 22179 13151 22185
rect 16206 22176 16212 22228
rect 16264 22216 16270 22228
rect 19337 22219 19395 22225
rect 19337 22216 19349 22219
rect 16264 22188 19349 22216
rect 16264 22176 16270 22188
rect 19337 22185 19349 22188
rect 19383 22185 19395 22219
rect 19337 22179 19395 22185
rect 20622 22176 20628 22228
rect 20680 22216 20686 22228
rect 21818 22216 21824 22228
rect 20680 22188 21824 22216
rect 20680 22176 20686 22188
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 22557 22219 22615 22225
rect 22557 22185 22569 22219
rect 22603 22216 22615 22219
rect 23198 22216 23204 22228
rect 22603 22188 23204 22216
rect 22603 22185 22615 22188
rect 22557 22179 22615 22185
rect 23198 22176 23204 22188
rect 23256 22176 23262 22228
rect 24578 22216 24584 22228
rect 23492 22188 24440 22216
rect 24539 22188 24584 22216
rect 16393 22151 16451 22157
rect 16393 22117 16405 22151
rect 16439 22148 16451 22151
rect 16666 22148 16672 22160
rect 16439 22120 16672 22148
rect 16439 22117 16451 22120
rect 16393 22111 16451 22117
rect 16666 22108 16672 22120
rect 16724 22108 16730 22160
rect 17497 22151 17555 22157
rect 17497 22117 17509 22151
rect 17543 22148 17555 22151
rect 20346 22148 20352 22160
rect 17543 22120 20352 22148
rect 17543 22117 17555 22120
rect 17497 22111 17555 22117
rect 20346 22108 20352 22120
rect 20404 22108 20410 22160
rect 20898 22148 20904 22160
rect 20456 22120 20904 22148
rect 8389 22083 8447 22089
rect 8389 22080 8401 22083
rect 7432 22052 8401 22080
rect 7432 22040 7438 22052
rect 8389 22049 8401 22052
rect 8435 22049 8447 22083
rect 8389 22043 8447 22049
rect 9401 22083 9459 22089
rect 9401 22049 9413 22083
rect 9447 22049 9459 22083
rect 13354 22080 13360 22092
rect 13315 22052 13360 22080
rect 9401 22043 9459 22049
rect 13354 22040 13360 22052
rect 13412 22040 13418 22092
rect 15841 22083 15899 22089
rect 15841 22049 15853 22083
rect 15887 22080 15899 22083
rect 16022 22080 16028 22092
rect 15887 22052 16028 22080
rect 15887 22049 15899 22052
rect 15841 22043 15899 22049
rect 16022 22040 16028 22052
rect 16080 22040 16086 22092
rect 17034 22080 17040 22092
rect 16995 22052 17040 22080
rect 17034 22040 17040 22052
rect 17092 22080 17098 22092
rect 17402 22080 17408 22092
rect 17092 22052 17408 22080
rect 17092 22040 17098 22052
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 18414 22080 18420 22092
rect 18375 22052 18420 22080
rect 18414 22040 18420 22052
rect 18472 22040 18478 22092
rect 18598 22080 18604 22092
rect 18559 22052 18604 22080
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 19705 22083 19763 22089
rect 19705 22049 19717 22083
rect 19751 22080 19763 22083
rect 20456 22080 20484 22120
rect 20898 22108 20904 22120
rect 20956 22108 20962 22160
rect 22925 22151 22983 22157
rect 22925 22117 22937 22151
rect 22971 22148 22983 22151
rect 23492 22148 23520 22188
rect 22971 22120 23520 22148
rect 22971 22117 22983 22120
rect 22925 22111 22983 22117
rect 23566 22108 23572 22160
rect 23624 22148 23630 22160
rect 24026 22148 24032 22160
rect 23624 22120 24032 22148
rect 23624 22108 23630 22120
rect 24026 22108 24032 22120
rect 24084 22108 24090 22160
rect 24412 22148 24440 22188
rect 24578 22176 24584 22188
rect 24636 22176 24642 22228
rect 28534 22176 28540 22228
rect 28592 22216 28598 22228
rect 28905 22219 28963 22225
rect 28905 22216 28917 22219
rect 28592 22188 28917 22216
rect 28592 22176 28598 22188
rect 28905 22185 28917 22188
rect 28951 22185 28963 22219
rect 28905 22179 28963 22185
rect 29917 22219 29975 22225
rect 29917 22185 29929 22219
rect 29963 22216 29975 22219
rect 30098 22216 30104 22228
rect 29963 22188 30104 22216
rect 29963 22185 29975 22188
rect 29917 22179 29975 22185
rect 30098 22176 30104 22188
rect 30156 22176 30162 22228
rect 36988 22219 37046 22225
rect 36988 22185 37000 22219
rect 37034 22216 37046 22219
rect 39206 22216 39212 22228
rect 37034 22188 39212 22216
rect 37034 22185 37046 22188
rect 36988 22179 37046 22185
rect 39206 22176 39212 22188
rect 39264 22176 39270 22228
rect 45646 22176 45652 22228
rect 45704 22216 45710 22228
rect 49142 22216 49148 22228
rect 45704 22188 49148 22216
rect 45704 22176 45710 22188
rect 49142 22176 49148 22188
rect 49200 22176 49206 22228
rect 49602 22216 49608 22228
rect 49563 22188 49608 22216
rect 49602 22176 49608 22188
rect 49660 22176 49666 22228
rect 51169 22219 51227 22225
rect 51169 22185 51181 22219
rect 51215 22216 51227 22219
rect 51978 22219 52036 22225
rect 51978 22216 51990 22219
rect 51215 22188 51990 22216
rect 51215 22185 51227 22188
rect 51169 22179 51227 22185
rect 51978 22185 51990 22188
rect 52024 22185 52036 22219
rect 51978 22179 52036 22185
rect 25682 22148 25688 22160
rect 24412 22120 25688 22148
rect 25682 22108 25688 22120
rect 25740 22108 25746 22160
rect 27798 22148 27804 22160
rect 27759 22120 27804 22148
rect 27798 22108 27804 22120
rect 27856 22108 27862 22160
rect 27893 22151 27951 22157
rect 27893 22117 27905 22151
rect 27939 22148 27951 22151
rect 28810 22148 28816 22160
rect 27939 22120 28816 22148
rect 27939 22117 27951 22120
rect 27893 22111 27951 22117
rect 28810 22108 28816 22120
rect 28868 22108 28874 22160
rect 40770 22108 40776 22160
rect 40828 22148 40834 22160
rect 44910 22148 44916 22160
rect 40828 22120 44916 22148
rect 40828 22108 40834 22120
rect 44910 22108 44916 22120
rect 44968 22108 44974 22160
rect 49620 22148 49648 22176
rect 48700 22120 49648 22148
rect 19751 22052 20484 22080
rect 19751 22049 19763 22052
rect 19705 22043 19763 22049
rect 21082 22040 21088 22092
rect 21140 22080 21146 22092
rect 21140 22052 23428 22080
rect 21140 22040 21146 22052
rect 1949 22015 2007 22021
rect 1949 21981 1961 22015
rect 1995 22012 2007 22015
rect 2866 22012 2872 22024
rect 1995 21984 2872 22012
rect 1995 21981 2007 21984
rect 1949 21975 2007 21981
rect 2866 21972 2872 21984
rect 2924 21972 2930 22024
rect 3234 22012 3240 22024
rect 3195 21984 3240 22012
rect 3234 21972 3240 21984
rect 3292 22012 3298 22024
rect 3789 22015 3847 22021
rect 3789 22012 3801 22015
rect 3292 21984 3801 22012
rect 3292 21972 3298 21984
rect 3789 21981 3801 21984
rect 3835 21981 3847 22015
rect 16298 22012 16304 22024
rect 16211 21984 16304 22012
rect 3789 21975 3847 21981
rect 16298 21972 16304 21984
rect 16356 22012 16362 22024
rect 16356 21984 16436 22012
rect 16356 21972 16362 21984
rect 6178 21944 6184 21956
rect 6139 21916 6184 21944
rect 6178 21904 6184 21916
rect 6236 21904 6242 21956
rect 7650 21904 7656 21956
rect 7708 21904 7714 21956
rect 8018 21904 8024 21956
rect 8076 21944 8082 21956
rect 8113 21947 8171 21953
rect 8113 21944 8125 21947
rect 8076 21916 8125 21944
rect 8076 21904 8082 21916
rect 8113 21913 8125 21916
rect 8159 21913 8171 21947
rect 9674 21944 9680 21956
rect 9635 21916 9680 21944
rect 8113 21907 8171 21913
rect 9674 21904 9680 21916
rect 9732 21904 9738 21956
rect 10134 21904 10140 21956
rect 10192 21904 10198 21956
rect 12434 21904 12440 21956
rect 12492 21904 12498 21956
rect 13722 21904 13728 21956
rect 13780 21944 13786 21956
rect 13780 21916 14320 21944
rect 13780 21904 13786 21916
rect 2866 21836 2872 21888
rect 2924 21876 2930 21888
rect 3145 21879 3203 21885
rect 3145 21876 3157 21879
rect 2924 21848 3157 21876
rect 2924 21836 2930 21848
rect 3145 21845 3157 21848
rect 3191 21845 3203 21879
rect 3145 21839 3203 21845
rect 3694 21836 3700 21888
rect 3752 21876 3758 21888
rect 6641 21879 6699 21885
rect 6641 21876 6653 21879
rect 3752 21848 6653 21876
rect 3752 21836 3758 21848
rect 6641 21845 6653 21848
rect 6687 21845 6699 21879
rect 6641 21839 6699 21845
rect 6730 21836 6736 21888
rect 6788 21876 6794 21888
rect 8938 21876 8944 21888
rect 6788 21848 8944 21876
rect 6788 21836 6794 21848
rect 8938 21836 8944 21848
rect 8996 21836 9002 21888
rect 11146 21876 11152 21888
rect 11107 21848 11152 21876
rect 11146 21836 11152 21848
rect 11204 21836 11210 21888
rect 11606 21876 11612 21888
rect 11567 21848 11612 21876
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 14090 21876 14096 21888
rect 14051 21848 14096 21876
rect 14090 21836 14096 21848
rect 14148 21836 14154 21888
rect 14292 21876 14320 21916
rect 15010 21904 15016 21956
rect 15068 21904 15074 21956
rect 15565 21947 15623 21953
rect 15565 21913 15577 21947
rect 15611 21944 15623 21947
rect 15838 21944 15844 21956
rect 15611 21916 15844 21944
rect 15611 21913 15623 21916
rect 15565 21907 15623 21913
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 16408 21944 16436 21984
rect 16482 21972 16488 22024
rect 16540 22012 16546 22024
rect 17129 22015 17187 22021
rect 17129 22012 17141 22015
rect 16540 21984 17141 22012
rect 16540 21972 16546 21984
rect 17129 21981 17141 21984
rect 17175 21981 17187 22015
rect 19334 22012 19340 22024
rect 17129 21975 17187 21981
rect 17236 21984 19340 22012
rect 17236 21944 17264 21984
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 19610 22012 19616 22024
rect 19571 21984 19616 22012
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 20349 22015 20407 22021
rect 20349 21981 20361 22015
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 22012 20591 22015
rect 20622 22012 20628 22024
rect 20579 21984 20628 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 16408 21916 17264 21944
rect 19150 21904 19156 21956
rect 19208 21944 19214 21956
rect 20364 21944 20392 21975
rect 20622 21972 20628 21984
rect 20680 21972 20686 22024
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 22012 21235 22015
rect 22462 22012 22468 22024
rect 21223 21984 21772 22012
rect 22423 21984 22468 22012
rect 21223 21981 21235 21984
rect 21177 21975 21235 21981
rect 19208 21916 20392 21944
rect 19208 21904 19214 21916
rect 17957 21879 18015 21885
rect 17957 21876 17969 21879
rect 14292 21848 17969 21876
rect 17957 21845 17969 21848
rect 18003 21845 18015 21879
rect 17957 21839 18015 21845
rect 18325 21879 18383 21885
rect 18325 21845 18337 21879
rect 18371 21876 18383 21879
rect 20162 21876 20168 21888
rect 18371 21848 20168 21876
rect 18371 21845 18383 21848
rect 18325 21839 18383 21845
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 20364 21876 20392 21916
rect 20441 21947 20499 21953
rect 20441 21913 20453 21947
rect 20487 21944 20499 21947
rect 21008 21944 21036 21975
rect 21637 21947 21695 21953
rect 21637 21944 21649 21947
rect 20487 21916 21649 21944
rect 20487 21913 20499 21916
rect 20441 21907 20499 21913
rect 21637 21913 21649 21916
rect 21683 21913 21695 21947
rect 21637 21907 21695 21913
rect 20990 21876 20996 21888
rect 20364 21848 20996 21876
rect 20990 21836 20996 21848
rect 21048 21836 21054 21888
rect 21082 21836 21088 21888
rect 21140 21876 21146 21888
rect 21744 21876 21772 21984
rect 22462 21972 22468 21984
rect 22520 21972 22526 22024
rect 22738 22012 22744 22024
rect 22699 21984 22744 22012
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 23400 22021 23428 22052
rect 25774 22040 25780 22092
rect 25832 22080 25838 22092
rect 26256 22083 26314 22089
rect 26256 22080 26268 22083
rect 25832 22052 26268 22080
rect 25832 22040 25838 22052
rect 26256 22049 26268 22052
rect 26302 22049 26314 22083
rect 29730 22080 29736 22092
rect 26256 22043 26314 22049
rect 27080 22052 29736 22080
rect 23385 22015 23443 22021
rect 23385 21981 23397 22015
rect 23431 21981 23443 22015
rect 23385 21975 23443 21981
rect 24394 21972 24400 22024
rect 24452 22012 24458 22024
rect 24489 22015 24547 22021
rect 24489 22012 24501 22015
rect 24452 21984 24501 22012
rect 24452 21972 24458 21984
rect 24489 21981 24501 21984
rect 24535 21981 24547 22015
rect 24489 21975 24547 21981
rect 24673 22015 24731 22021
rect 24673 21981 24685 22015
rect 24719 22012 24731 22015
rect 24946 22012 24952 22024
rect 24719 21984 24952 22012
rect 24719 21981 24731 21984
rect 24673 21975 24731 21981
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 25590 22012 25596 22024
rect 25551 21984 25596 22012
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 26050 22012 26056 22024
rect 26011 21984 26056 22012
rect 26050 21972 26056 21984
rect 26108 21972 26114 22024
rect 26510 22012 26516 22024
rect 26206 21984 26516 22012
rect 21818 21904 21824 21956
rect 21876 21944 21882 21956
rect 22005 21947 22063 21953
rect 21876 21916 21921 21944
rect 21876 21904 21882 21916
rect 22005 21913 22017 21947
rect 22051 21944 22063 21947
rect 23842 21944 23848 21956
rect 22051 21916 23848 21944
rect 22051 21913 22063 21916
rect 22005 21907 22063 21913
rect 23842 21904 23848 21916
rect 23900 21904 23906 21956
rect 24210 21904 24216 21956
rect 24268 21944 24274 21956
rect 25958 21944 25964 21956
rect 24268 21916 25964 21944
rect 24268 21904 24274 21916
rect 25958 21904 25964 21916
rect 26016 21944 26022 21956
rect 26206 21944 26234 21984
rect 26510 21972 26516 21984
rect 26568 22012 26574 22024
rect 27080 22021 27108 22052
rect 29730 22040 29736 22052
rect 29788 22040 29794 22092
rect 31570 22080 31576 22092
rect 31531 22052 31576 22080
rect 31570 22040 31576 22052
rect 31628 22040 31634 22092
rect 33870 22040 33876 22092
rect 33928 22080 33934 22092
rect 34057 22083 34115 22089
rect 34057 22080 34069 22083
rect 33928 22052 34069 22080
rect 33928 22040 33934 22052
rect 34057 22049 34069 22052
rect 34103 22049 34115 22083
rect 34057 22043 34115 22049
rect 38473 22083 38531 22089
rect 38473 22049 38485 22083
rect 38519 22049 38531 22083
rect 45278 22080 45284 22092
rect 38473 22043 38531 22049
rect 43824 22052 45284 22080
rect 26881 22015 26939 22021
rect 26881 22012 26893 22015
rect 26568 21984 26893 22012
rect 26568 21972 26574 21984
rect 26881 21981 26893 21984
rect 26927 21981 26939 22015
rect 26881 21975 26939 21981
rect 27065 22015 27123 22021
rect 27065 21981 27077 22015
rect 27111 21981 27123 22015
rect 27065 21975 27123 21981
rect 27154 21972 27160 22024
rect 27212 22012 27218 22024
rect 27709 22015 27767 22021
rect 27709 22012 27721 22015
rect 27212 21984 27721 22012
rect 27212 21972 27218 21984
rect 27709 21981 27721 21984
rect 27755 21981 27767 22015
rect 27709 21975 27767 21981
rect 26016 21916 26234 21944
rect 26329 21947 26387 21953
rect 26016 21904 26022 21916
rect 26329 21913 26341 21947
rect 26375 21944 26387 21947
rect 27525 21947 27583 21953
rect 27525 21944 27537 21947
rect 26375 21916 27537 21944
rect 26375 21913 26387 21916
rect 26329 21907 26387 21913
rect 27525 21913 27537 21916
rect 27571 21913 27583 21947
rect 27525 21907 27583 21913
rect 24486 21876 24492 21888
rect 21140 21848 21185 21876
rect 21744 21848 24492 21876
rect 21140 21836 21146 21848
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 24854 21876 24860 21888
rect 24815 21848 24860 21876
rect 24854 21836 24860 21848
rect 24912 21836 24918 21888
rect 25498 21876 25504 21888
rect 25459 21848 25504 21876
rect 25498 21836 25504 21848
rect 25556 21836 25562 21888
rect 26142 21876 26148 21888
rect 26103 21848 26148 21876
rect 26142 21836 26148 21848
rect 26200 21836 26206 21888
rect 26973 21879 27031 21885
rect 26973 21845 26985 21879
rect 27019 21876 27031 21879
rect 27338 21876 27344 21888
rect 27019 21848 27344 21876
rect 27019 21845 27031 21848
rect 26973 21839 27031 21845
rect 27338 21836 27344 21848
rect 27396 21836 27402 21888
rect 27724 21876 27752 21975
rect 27982 21972 27988 22024
rect 28040 22012 28046 22024
rect 28169 22015 28227 22021
rect 28040 21984 28085 22012
rect 28040 21972 28046 21984
rect 28169 21981 28181 22015
rect 28215 21981 28227 22015
rect 28169 21975 28227 21981
rect 28184 21944 28212 21975
rect 28258 21972 28264 22024
rect 28316 22012 28322 22024
rect 28813 22015 28871 22021
rect 28813 22012 28825 22015
rect 28316 21984 28825 22012
rect 28316 21972 28322 21984
rect 28813 21981 28825 21984
rect 28859 21981 28871 22015
rect 28994 22012 29000 22024
rect 28955 21984 29000 22012
rect 28813 21975 28871 21981
rect 28994 21972 29000 21984
rect 29052 21972 29058 22024
rect 30009 22015 30067 22021
rect 30009 21981 30021 22015
rect 30055 21981 30067 22015
rect 30466 22012 30472 22024
rect 30427 21984 30472 22012
rect 30009 21975 30067 21981
rect 28350 21944 28356 21956
rect 28184 21916 28356 21944
rect 28350 21904 28356 21916
rect 28408 21904 28414 21956
rect 30024 21944 30052 21975
rect 30466 21972 30472 21984
rect 30524 21972 30530 22024
rect 31481 22015 31539 22021
rect 31481 21981 31493 22015
rect 31527 21981 31539 22015
rect 34146 22012 34152 22024
rect 34059 21984 34152 22012
rect 31481 21975 31539 21981
rect 31294 21944 31300 21956
rect 30024 21916 31300 21944
rect 31294 21904 31300 21916
rect 31352 21944 31358 21956
rect 31496 21944 31524 21975
rect 34146 21972 34152 21984
rect 34204 22012 34210 22024
rect 35253 22015 35311 22021
rect 35253 22012 35265 22015
rect 34204 21984 35265 22012
rect 34204 21972 34210 21984
rect 35253 21981 35265 21984
rect 35299 21981 35311 22015
rect 35253 21975 35311 21981
rect 35621 22015 35679 22021
rect 35621 21981 35633 22015
rect 35667 22012 35679 22015
rect 35894 22012 35900 22024
rect 35667 21984 35900 22012
rect 35667 21981 35679 21984
rect 35621 21975 35679 21981
rect 35894 21972 35900 21984
rect 35952 21972 35958 22024
rect 36722 22012 36728 22024
rect 36683 21984 36728 22012
rect 36722 21972 36728 21984
rect 36780 21972 36786 22024
rect 38488 22012 38516 22043
rect 39209 22015 39267 22021
rect 39209 22012 39221 22015
rect 38488 21984 39221 22012
rect 39209 21981 39221 21984
rect 39255 22012 39267 22015
rect 39298 22012 39304 22024
rect 39255 21984 39304 22012
rect 39255 21981 39267 21984
rect 39209 21975 39267 21981
rect 39298 21972 39304 21984
rect 39356 21972 39362 22024
rect 40034 22012 40040 22024
rect 39995 21984 40040 22012
rect 40034 21972 40040 21984
rect 40092 21972 40098 22024
rect 43438 21972 43444 22024
rect 43496 22012 43502 22024
rect 43625 22015 43683 22021
rect 43625 22012 43637 22015
rect 43496 21984 43637 22012
rect 43496 21972 43502 21984
rect 43625 21981 43637 21984
rect 43671 21981 43683 22015
rect 43625 21975 43683 21981
rect 31352 21916 31524 21944
rect 31352 21904 31358 21916
rect 37734 21904 37740 21956
rect 37792 21904 37798 21956
rect 29454 21876 29460 21888
rect 27724 21848 29460 21876
rect 29454 21836 29460 21848
rect 29512 21836 29518 21888
rect 30558 21876 30564 21888
rect 30519 21848 30564 21876
rect 30558 21836 30564 21848
rect 30616 21836 30622 21888
rect 32306 21876 32312 21888
rect 32267 21848 32312 21876
rect 32306 21836 32312 21848
rect 32364 21836 32370 21888
rect 36265 21879 36323 21885
rect 36265 21845 36277 21879
rect 36311 21876 36323 21879
rect 36906 21876 36912 21888
rect 36311 21848 36912 21876
rect 36311 21845 36323 21848
rect 36265 21839 36323 21845
rect 36906 21836 36912 21848
rect 36964 21836 36970 21888
rect 38562 21836 38568 21888
rect 38620 21876 38626 21888
rect 39025 21879 39083 21885
rect 39025 21876 39037 21879
rect 38620 21848 39037 21876
rect 38620 21836 38626 21848
rect 39025 21845 39037 21848
rect 39071 21845 39083 21879
rect 39025 21839 39083 21845
rect 39482 21836 39488 21888
rect 39540 21876 39546 21888
rect 43824 21885 43852 22052
rect 45278 22040 45284 22052
rect 45336 22040 45342 22092
rect 45465 22083 45523 22089
rect 45465 22049 45477 22083
rect 45511 22080 45523 22083
rect 47210 22080 47216 22092
rect 45511 22052 47216 22080
rect 45511 22049 45523 22052
rect 45465 22043 45523 22049
rect 47210 22040 47216 22052
rect 47268 22040 47274 22092
rect 48314 22080 48320 22092
rect 48275 22052 48320 22080
rect 48314 22040 48320 22052
rect 48372 22040 48378 22092
rect 44082 21972 44088 22024
rect 44140 22012 44146 22024
rect 44269 22015 44327 22021
rect 44269 22012 44281 22015
rect 44140 21984 44281 22012
rect 44140 21972 44146 21984
rect 44269 21981 44281 21984
rect 44315 21981 44327 22015
rect 45370 22012 45376 22024
rect 45331 21984 45376 22012
rect 44269 21975 44327 21981
rect 45370 21972 45376 21984
rect 45428 21972 45434 22024
rect 46198 21972 46204 22024
rect 46256 22012 46262 22024
rect 47397 22015 47455 22021
rect 47397 22012 47409 22015
rect 46256 21984 47409 22012
rect 46256 21972 46262 21984
rect 47397 21981 47409 21984
rect 47443 21981 47455 22015
rect 47397 21975 47455 21981
rect 47762 21972 47768 22024
rect 47820 22012 47826 22024
rect 48225 22015 48283 22021
rect 48225 22012 48237 22015
rect 47820 21984 48237 22012
rect 47820 21972 47826 21984
rect 48225 21981 48237 21984
rect 48271 22012 48283 22015
rect 48700 22012 48728 22120
rect 49513 22083 49571 22089
rect 49513 22049 49525 22083
rect 49559 22080 49571 22083
rect 49559 22052 50568 22080
rect 49559 22049 49571 22052
rect 49513 22043 49571 22049
rect 48271 21984 48728 22012
rect 49605 22015 49663 22021
rect 48271 21981 48283 21984
rect 48225 21975 48283 21981
rect 49605 21981 49617 22015
rect 49651 22012 49663 22015
rect 50154 22012 50160 22024
rect 49651 21984 50160 22012
rect 49651 21981 49663 21984
rect 49605 21975 49663 21981
rect 50154 21972 50160 21984
rect 50212 21972 50218 22024
rect 50540 22012 50568 22052
rect 50614 22040 50620 22092
rect 50672 22080 50678 22092
rect 50801 22083 50859 22089
rect 50801 22080 50813 22083
rect 50672 22052 50813 22080
rect 50672 22040 50678 22052
rect 50801 22049 50813 22052
rect 50847 22049 50859 22083
rect 53469 22083 53527 22089
rect 53469 22080 53481 22083
rect 50801 22043 50859 22049
rect 51046 22052 53481 22080
rect 50706 22012 50712 22024
rect 50540 21984 50712 22012
rect 50706 21972 50712 21984
rect 50764 22012 50770 22024
rect 50893 22015 50951 22021
rect 50893 22012 50905 22015
rect 50764 21984 50905 22012
rect 50764 21972 50770 21984
rect 50893 21981 50905 21984
rect 50939 22012 50951 22015
rect 51046 22012 51074 22052
rect 53469 22049 53481 22052
rect 53515 22049 53527 22083
rect 53469 22043 53527 22049
rect 50939 21984 51074 22012
rect 51721 22015 51779 22021
rect 50939 21981 50951 21984
rect 50893 21975 50951 21981
rect 51721 21981 51733 22015
rect 51767 21981 51779 22015
rect 51721 21975 51779 21981
rect 45278 21904 45284 21956
rect 45336 21944 45342 21956
rect 48406 21944 48412 21956
rect 45336 21916 48412 21944
rect 45336 21904 45342 21916
rect 48406 21904 48412 21916
rect 48464 21944 48470 21956
rect 51736 21944 51764 21975
rect 55122 21972 55128 22024
rect 55180 22012 55186 22024
rect 55401 22015 55459 22021
rect 55401 22012 55413 22015
rect 55180 21984 55413 22012
rect 55180 21972 55186 21984
rect 55401 21981 55413 21984
rect 55447 21981 55459 22015
rect 55401 21975 55459 21981
rect 51902 21944 51908 21956
rect 48464 21916 51908 21944
rect 48464 21904 48470 21916
rect 51902 21904 51908 21916
rect 51960 21904 51966 21956
rect 52380 21916 52486 21944
rect 52380 21888 52408 21916
rect 39945 21879 40003 21885
rect 39945 21876 39957 21879
rect 39540 21848 39957 21876
rect 39540 21836 39546 21848
rect 39945 21845 39957 21848
rect 39991 21845 40003 21879
rect 39945 21839 40003 21845
rect 43809 21879 43867 21885
rect 43809 21845 43821 21879
rect 43855 21845 43867 21879
rect 43809 21839 43867 21845
rect 44174 21836 44180 21888
rect 44232 21876 44238 21888
rect 44453 21879 44511 21885
rect 44453 21876 44465 21879
rect 44232 21848 44465 21876
rect 44232 21836 44238 21848
rect 44453 21845 44465 21848
rect 44499 21845 44511 21879
rect 45002 21876 45008 21888
rect 44963 21848 45008 21876
rect 44453 21839 44511 21845
rect 45002 21836 45008 21848
rect 45060 21836 45066 21888
rect 45738 21836 45744 21888
rect 45796 21876 45802 21888
rect 46017 21879 46075 21885
rect 46017 21876 46029 21879
rect 45796 21848 46029 21876
rect 45796 21836 45802 21848
rect 46017 21845 46029 21848
rect 46063 21876 46075 21879
rect 46566 21876 46572 21888
rect 46063 21848 46572 21876
rect 46063 21845 46075 21848
rect 46017 21839 46075 21845
rect 46566 21836 46572 21848
rect 46624 21836 46630 21888
rect 47578 21876 47584 21888
rect 47539 21848 47584 21876
rect 47578 21836 47584 21848
rect 47636 21836 47642 21888
rect 48590 21876 48596 21888
rect 48551 21848 48596 21876
rect 48590 21836 48596 21848
rect 48648 21836 48654 21888
rect 49234 21876 49240 21888
rect 49195 21848 49240 21876
rect 49234 21836 49240 21848
rect 49292 21836 49298 21888
rect 49970 21836 49976 21888
rect 50028 21876 50034 21888
rect 50157 21879 50215 21885
rect 50157 21876 50169 21879
rect 50028 21848 50169 21876
rect 50028 21836 50034 21848
rect 50157 21845 50169 21848
rect 50203 21845 50215 21879
rect 50157 21839 50215 21845
rect 52362 21836 52368 21888
rect 52420 21836 52426 21888
rect 55582 21876 55588 21888
rect 55543 21848 55588 21876
rect 55582 21836 55588 21848
rect 55640 21836 55646 21888
rect 1104 21786 58880 21808
rect 1104 21734 15398 21786
rect 15450 21734 15462 21786
rect 15514 21734 15526 21786
rect 15578 21734 15590 21786
rect 15642 21734 15654 21786
rect 15706 21734 29846 21786
rect 29898 21734 29910 21786
rect 29962 21734 29974 21786
rect 30026 21734 30038 21786
rect 30090 21734 30102 21786
rect 30154 21734 44294 21786
rect 44346 21734 44358 21786
rect 44410 21734 44422 21786
rect 44474 21734 44486 21786
rect 44538 21734 44550 21786
rect 44602 21734 58880 21786
rect 1104 21712 58880 21734
rect 1857 21675 1915 21681
rect 1857 21641 1869 21675
rect 1903 21672 1915 21675
rect 3970 21672 3976 21684
rect 1903 21644 3976 21672
rect 1903 21641 1915 21644
rect 1857 21635 1915 21641
rect 3970 21632 3976 21644
rect 4028 21632 4034 21684
rect 4065 21675 4123 21681
rect 4065 21641 4077 21675
rect 4111 21672 4123 21675
rect 4111 21644 6132 21672
rect 4111 21641 4123 21644
rect 4065 21635 4123 21641
rect 2866 21564 2872 21616
rect 2924 21564 2930 21616
rect 5442 21604 5448 21616
rect 5106 21576 5448 21604
rect 5442 21564 5448 21576
rect 5500 21564 5506 21616
rect 5537 21607 5595 21613
rect 5537 21573 5549 21607
rect 5583 21604 5595 21607
rect 5902 21604 5908 21616
rect 5583 21576 5908 21604
rect 5583 21573 5595 21576
rect 5537 21567 5595 21573
rect 5902 21564 5908 21576
rect 5960 21564 5966 21616
rect 6104 21604 6132 21644
rect 6178 21632 6184 21684
rect 6236 21672 6242 21684
rect 11790 21672 11796 21684
rect 6236 21644 8708 21672
rect 11751 21644 11796 21672
rect 6236 21632 6242 21644
rect 6730 21604 6736 21616
rect 6104 21576 6736 21604
rect 6730 21564 6736 21576
rect 6788 21564 6794 21616
rect 7098 21564 7104 21616
rect 7156 21564 7162 21616
rect 8680 21613 8708 21644
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 13170 21632 13176 21684
rect 13228 21672 13234 21684
rect 14737 21675 14795 21681
rect 14737 21672 14749 21675
rect 13228 21644 14749 21672
rect 13228 21632 13234 21644
rect 14737 21641 14749 21644
rect 14783 21641 14795 21675
rect 14737 21635 14795 21641
rect 17954 21632 17960 21684
rect 18012 21672 18018 21684
rect 18417 21675 18475 21681
rect 18417 21672 18429 21675
rect 18012 21644 18429 21672
rect 18012 21632 18018 21644
rect 18417 21641 18429 21644
rect 18463 21641 18475 21675
rect 18417 21635 18475 21641
rect 20162 21632 20168 21684
rect 20220 21672 20226 21684
rect 21082 21672 21088 21684
rect 20220 21644 21088 21672
rect 20220 21632 20226 21644
rect 21082 21632 21088 21644
rect 21140 21632 21146 21684
rect 24946 21672 24952 21684
rect 22066 21644 24952 21672
rect 8665 21607 8723 21613
rect 8665 21573 8677 21607
rect 8711 21604 8723 21607
rect 9398 21604 9404 21616
rect 8711 21576 9404 21604
rect 8711 21573 8723 21576
rect 8665 21567 8723 21573
rect 9398 21564 9404 21576
rect 9456 21564 9462 21616
rect 10965 21607 11023 21613
rect 10965 21573 10977 21607
rect 11011 21604 11023 21607
rect 16298 21604 16304 21616
rect 11011 21576 16304 21604
rect 11011 21573 11023 21576
rect 10965 21567 11023 21573
rect 5810 21496 5816 21548
rect 5868 21536 5874 21548
rect 10410 21536 10416 21548
rect 5868 21508 5913 21536
rect 10371 21508 10416 21536
rect 5868 21496 5874 21508
rect 10410 21496 10416 21508
rect 10468 21496 10474 21548
rect 3326 21468 3332 21480
rect 3287 21440 3332 21468
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 3602 21468 3608 21480
rect 3563 21440 3608 21468
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 4338 21428 4344 21480
rect 4396 21468 4402 21480
rect 6365 21471 6423 21477
rect 6365 21468 6377 21471
rect 4396 21440 6377 21468
rect 4396 21428 4402 21440
rect 6365 21437 6377 21440
rect 6411 21437 6423 21471
rect 6641 21471 6699 21477
rect 6641 21468 6653 21471
rect 6365 21431 6423 21437
rect 6472 21440 6653 21468
rect 5074 21292 5080 21344
rect 5132 21332 5138 21344
rect 6472 21332 6500 21440
rect 6641 21437 6653 21440
rect 6687 21437 6699 21471
rect 6641 21431 6699 21437
rect 6730 21428 6736 21480
rect 6788 21468 6794 21480
rect 10980 21468 11008 21567
rect 16298 21564 16304 21576
rect 16356 21564 16362 21616
rect 17126 21604 17132 21616
rect 17087 21576 17132 21604
rect 17126 21564 17132 21576
rect 17184 21564 17190 21616
rect 19610 21604 19616 21616
rect 18524 21576 19616 21604
rect 11698 21536 11704 21548
rect 11659 21508 11704 21536
rect 11698 21496 11704 21508
rect 11756 21496 11762 21548
rect 11790 21496 11796 21548
rect 11848 21536 11854 21548
rect 12345 21539 12403 21545
rect 12345 21536 12357 21539
rect 11848 21508 12357 21536
rect 11848 21496 11854 21508
rect 12345 21505 12357 21508
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 14921 21539 14979 21545
rect 14921 21505 14933 21539
rect 14967 21536 14979 21539
rect 15010 21536 15016 21548
rect 14967 21508 15016 21536
rect 14967 21505 14979 21508
rect 14921 21499 14979 21505
rect 15010 21496 15016 21508
rect 15068 21496 15074 21548
rect 15746 21536 15752 21548
rect 15707 21508 15752 21536
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 16390 21496 16396 21548
rect 16448 21536 16454 21548
rect 18524 21536 18552 21576
rect 18690 21536 18696 21548
rect 16448 21508 18552 21536
rect 18651 21508 18696 21536
rect 16448 21496 16454 21508
rect 18690 21496 18696 21508
rect 18748 21496 18754 21548
rect 19444 21545 19472 21576
rect 19610 21564 19616 21576
rect 19668 21564 19674 21616
rect 22066 21604 22094 21644
rect 24946 21632 24952 21644
rect 25004 21632 25010 21684
rect 25590 21632 25596 21684
rect 25648 21672 25654 21684
rect 27798 21672 27804 21684
rect 25648 21644 27804 21672
rect 25648 21632 25654 21644
rect 27798 21632 27804 21644
rect 27856 21632 27862 21684
rect 27890 21632 27896 21684
rect 27948 21672 27954 21684
rect 28077 21675 28135 21681
rect 28077 21672 28089 21675
rect 27948 21644 28089 21672
rect 27948 21632 27954 21644
rect 28077 21641 28089 21644
rect 28123 21641 28135 21675
rect 34241 21675 34299 21681
rect 34241 21672 34253 21675
rect 28077 21635 28135 21641
rect 33520 21644 34253 21672
rect 25498 21604 25504 21616
rect 20732 21576 22094 21604
rect 24794 21576 25504 21604
rect 19429 21539 19487 21545
rect 19429 21505 19441 21539
rect 19475 21505 19487 21539
rect 19429 21499 19487 21505
rect 20732 21480 20760 21576
rect 25498 21564 25504 21576
rect 25556 21564 25562 21616
rect 26050 21564 26056 21616
rect 26108 21564 26114 21616
rect 26878 21564 26884 21616
rect 26936 21604 26942 21616
rect 27522 21604 27528 21616
rect 26936 21576 27528 21604
rect 26936 21564 26942 21576
rect 27522 21564 27528 21576
rect 27580 21564 27586 21616
rect 27614 21564 27620 21616
rect 27672 21604 27678 21616
rect 28629 21607 28687 21613
rect 28629 21604 28641 21607
rect 27672 21576 28641 21604
rect 27672 21564 27678 21576
rect 28629 21573 28641 21576
rect 28675 21573 28687 21607
rect 30190 21604 30196 21616
rect 30151 21576 30196 21604
rect 28629 21567 28687 21573
rect 30190 21564 30196 21576
rect 30248 21564 30254 21616
rect 22278 21536 22284 21548
rect 22066 21508 22284 21536
rect 6788 21440 11008 21468
rect 6788 21428 6794 21440
rect 15286 21428 15292 21480
rect 15344 21468 15350 21480
rect 15381 21471 15439 21477
rect 15381 21468 15393 21471
rect 15344 21440 15393 21468
rect 15344 21428 15350 21440
rect 15381 21437 15393 21440
rect 15427 21437 15439 21471
rect 15381 21431 15439 21437
rect 15841 21471 15899 21477
rect 15841 21437 15853 21471
rect 15887 21468 15899 21471
rect 18322 21468 18328 21480
rect 15887 21440 18328 21468
rect 15887 21437 15899 21440
rect 15841 21431 15899 21437
rect 18322 21428 18328 21440
rect 18380 21428 18386 21480
rect 18417 21471 18475 21477
rect 18417 21437 18429 21471
rect 18463 21437 18475 21471
rect 18417 21431 18475 21437
rect 18601 21471 18659 21477
rect 18601 21437 18613 21471
rect 18647 21468 18659 21471
rect 19242 21468 19248 21480
rect 18647 21440 19248 21468
rect 18647 21437 18659 21440
rect 18601 21431 18659 21437
rect 10962 21360 10968 21412
rect 11020 21400 11026 21412
rect 17770 21400 17776 21412
rect 11020 21372 17776 21400
rect 11020 21360 11026 21372
rect 17770 21360 17776 21372
rect 17828 21400 17834 21412
rect 18432 21400 18460 21431
rect 19242 21428 19248 21440
rect 19300 21428 19306 21480
rect 19337 21471 19395 21477
rect 19337 21437 19349 21471
rect 19383 21437 19395 21471
rect 19794 21468 19800 21480
rect 19755 21440 19800 21468
rect 19337 21431 19395 21437
rect 17828 21372 18460 21400
rect 17828 21360 17834 21372
rect 19150 21360 19156 21412
rect 19208 21400 19214 21412
rect 19352 21400 19380 21431
rect 19794 21428 19800 21440
rect 19852 21468 19858 21480
rect 20257 21471 20315 21477
rect 20257 21468 20269 21471
rect 19852 21440 20269 21468
rect 19852 21428 19858 21440
rect 20257 21437 20269 21440
rect 20303 21437 20315 21471
rect 20257 21431 20315 21437
rect 20533 21471 20591 21477
rect 20533 21437 20545 21471
rect 20579 21468 20591 21471
rect 20714 21468 20720 21480
rect 20579 21440 20720 21468
rect 20579 21437 20591 21440
rect 20533 21431 20591 21437
rect 20714 21428 20720 21440
rect 20772 21428 20778 21480
rect 19208 21372 19380 21400
rect 19208 21360 19214 21372
rect 5132 21304 6500 21332
rect 5132 21292 5138 21304
rect 7190 21292 7196 21344
rect 7248 21332 7254 21344
rect 8113 21335 8171 21341
rect 8113 21332 8125 21335
rect 7248 21304 8125 21332
rect 7248 21292 7254 21304
rect 8113 21301 8125 21304
rect 8159 21301 8171 21335
rect 8113 21295 8171 21301
rect 12986 21292 12992 21344
rect 13044 21332 13050 21344
rect 13633 21335 13691 21341
rect 13633 21332 13645 21335
rect 13044 21304 13645 21332
rect 13044 21292 13050 21304
rect 13633 21301 13645 21304
rect 13679 21301 13691 21335
rect 13633 21295 13691 21301
rect 15746 21292 15752 21344
rect 15804 21332 15810 21344
rect 17402 21332 17408 21344
rect 15804 21304 17408 21332
rect 15804 21292 15810 21304
rect 17402 21292 17408 21304
rect 17460 21292 17466 21344
rect 19352 21332 19380 21372
rect 20346 21360 20352 21412
rect 20404 21400 20410 21412
rect 22066 21400 22094 21508
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 23290 21536 23296 21548
rect 23251 21508 23296 21536
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 24854 21496 24860 21548
rect 24912 21536 24918 21548
rect 25685 21539 25743 21545
rect 25685 21536 25697 21539
rect 24912 21508 25697 21536
rect 24912 21496 24918 21508
rect 25685 21505 25697 21508
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21536 25927 21539
rect 26068 21536 26096 21564
rect 26234 21536 26240 21548
rect 25915 21508 26096 21536
rect 26195 21508 26240 21536
rect 25915 21505 25927 21508
rect 25869 21499 25927 21505
rect 26234 21496 26240 21508
rect 26292 21496 26298 21548
rect 27154 21536 27160 21548
rect 27115 21508 27160 21536
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 27246 21496 27252 21548
rect 27304 21536 27310 21548
rect 27433 21539 27491 21545
rect 27433 21536 27445 21539
rect 27304 21508 27445 21536
rect 27304 21496 27310 21508
rect 27433 21505 27445 21508
rect 27479 21505 27491 21539
rect 27433 21499 27491 21505
rect 27890 21496 27896 21548
rect 27948 21536 27954 21548
rect 27985 21539 28043 21545
rect 27985 21536 27997 21539
rect 27948 21508 27997 21536
rect 27948 21496 27954 21508
rect 27985 21505 27997 21508
rect 28031 21505 28043 21539
rect 28166 21536 28172 21548
rect 28127 21508 28172 21536
rect 27985 21499 28043 21505
rect 28166 21496 28172 21508
rect 28224 21496 28230 21548
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21536 31263 21539
rect 31570 21536 31576 21548
rect 31251 21508 31576 21536
rect 31251 21505 31263 21508
rect 31205 21499 31263 21505
rect 31570 21496 31576 21508
rect 31628 21496 31634 21548
rect 32858 21536 32864 21548
rect 32819 21508 32864 21536
rect 32858 21496 32864 21508
rect 32916 21496 32922 21548
rect 33520 21545 33548 21644
rect 34241 21641 34253 21644
rect 34287 21672 34299 21675
rect 35434 21672 35440 21684
rect 34287 21644 35440 21672
rect 34287 21641 34299 21644
rect 34241 21635 34299 21641
rect 35434 21632 35440 21644
rect 35492 21632 35498 21684
rect 36262 21672 36268 21684
rect 36223 21644 36268 21672
rect 36262 21632 36268 21644
rect 36320 21632 36326 21684
rect 39758 21672 39764 21684
rect 39719 21644 39764 21672
rect 39758 21632 39764 21644
rect 39816 21672 39822 21684
rect 45370 21672 45376 21684
rect 39816 21644 40540 21672
rect 39816 21632 39822 21644
rect 35452 21604 35480 21632
rect 38289 21607 38347 21613
rect 35452 21576 37320 21604
rect 33505 21539 33563 21545
rect 33505 21505 33517 21539
rect 33551 21505 33563 21539
rect 33505 21499 33563 21505
rect 34425 21539 34483 21545
rect 34425 21505 34437 21539
rect 34471 21536 34483 21539
rect 34514 21536 34520 21548
rect 34471 21508 34520 21536
rect 34471 21505 34483 21508
rect 34425 21499 34483 21505
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 23658 21468 23664 21480
rect 23615 21440 23664 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 24946 21428 24952 21480
rect 25004 21428 25010 21480
rect 25961 21471 26019 21477
rect 25961 21437 25973 21471
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 26053 21471 26111 21477
rect 26053 21437 26065 21471
rect 26099 21468 26111 21471
rect 26973 21471 27031 21477
rect 26973 21468 26985 21471
rect 26099 21440 26985 21468
rect 26099 21437 26111 21440
rect 26053 21431 26111 21437
rect 26973 21437 26985 21440
rect 27019 21437 27031 21471
rect 26973 21431 27031 21437
rect 20404 21372 22094 21400
rect 24964 21400 24992 21428
rect 25866 21400 25872 21412
rect 24964 21372 25872 21400
rect 20404 21360 20410 21372
rect 25866 21360 25872 21372
rect 25924 21360 25930 21412
rect 25976 21400 26004 21431
rect 27062 21428 27068 21480
rect 27120 21468 27126 21480
rect 28074 21468 28080 21480
rect 27120 21440 28080 21468
rect 27120 21428 27126 21440
rect 26510 21400 26516 21412
rect 25976 21372 26516 21400
rect 26510 21360 26516 21372
rect 26568 21400 26574 21412
rect 26878 21400 26884 21412
rect 26568 21372 26884 21400
rect 26568 21360 26574 21372
rect 26878 21360 26884 21372
rect 26936 21360 26942 21412
rect 27264 21409 27292 21440
rect 28074 21428 28080 21440
rect 28132 21428 28138 21480
rect 30466 21428 30472 21480
rect 30524 21468 30530 21480
rect 33520 21468 33548 21499
rect 34514 21496 34520 21508
rect 34572 21536 34578 21548
rect 35437 21539 35495 21545
rect 35437 21536 35449 21539
rect 34572 21508 35449 21536
rect 34572 21496 34578 21508
rect 35437 21505 35449 21508
rect 35483 21536 35495 21539
rect 35618 21536 35624 21548
rect 35483 21508 35624 21536
rect 35483 21505 35495 21508
rect 35437 21499 35495 21505
rect 35618 21496 35624 21508
rect 35676 21536 35682 21548
rect 36449 21539 36507 21545
rect 36449 21536 36461 21539
rect 35676 21508 36461 21536
rect 35676 21496 35682 21508
rect 36449 21505 36461 21508
rect 36495 21536 36507 21539
rect 36998 21536 37004 21548
rect 36495 21508 37004 21536
rect 36495 21505 36507 21508
rect 36449 21499 36507 21505
rect 36998 21496 37004 21508
rect 37056 21496 37062 21548
rect 37292 21545 37320 21576
rect 38289 21573 38301 21607
rect 38335 21604 38347 21607
rect 38562 21604 38568 21616
rect 38335 21576 38568 21604
rect 38335 21573 38347 21576
rect 38289 21567 38347 21573
rect 38562 21564 38568 21576
rect 38620 21564 38626 21616
rect 40313 21607 40371 21613
rect 40313 21604 40325 21607
rect 39514 21576 40325 21604
rect 40313 21573 40325 21576
rect 40359 21573 40371 21607
rect 40313 21567 40371 21573
rect 37277 21539 37335 21545
rect 37277 21505 37289 21539
rect 37323 21505 37335 21539
rect 38010 21536 38016 21548
rect 37971 21508 38016 21536
rect 37277 21499 37335 21505
rect 38010 21496 38016 21508
rect 38068 21496 38074 21548
rect 40402 21536 40408 21548
rect 40363 21508 40408 21536
rect 40402 21496 40408 21508
rect 40460 21496 40466 21548
rect 40512 21536 40540 21644
rect 44284 21644 45376 21672
rect 44284 21545 44312 21644
rect 45370 21632 45376 21644
rect 45428 21672 45434 21684
rect 46523 21675 46581 21681
rect 46523 21672 46535 21675
rect 45428 21644 46535 21672
rect 45428 21632 45434 21644
rect 46523 21641 46535 21644
rect 46569 21641 46581 21675
rect 46523 21635 46581 21641
rect 47486 21632 47492 21684
rect 47544 21672 47550 21684
rect 47765 21675 47823 21681
rect 47765 21672 47777 21675
rect 47544 21644 47777 21672
rect 47544 21632 47550 21644
rect 47765 21641 47777 21644
rect 47811 21641 47823 21675
rect 49510 21672 49516 21684
rect 47765 21635 47823 21641
rect 48516 21644 49516 21672
rect 45646 21564 45652 21616
rect 45704 21564 45710 21616
rect 48516 21604 48544 21644
rect 49510 21632 49516 21644
rect 49568 21632 49574 21684
rect 49602 21632 49608 21684
rect 49660 21672 49666 21684
rect 50157 21675 50215 21681
rect 50157 21672 50169 21675
rect 49660 21644 50169 21672
rect 49660 21632 49666 21644
rect 50157 21641 50169 21644
rect 50203 21641 50215 21675
rect 50157 21635 50215 21641
rect 47688 21576 48544 21604
rect 47688 21548 47716 21576
rect 48590 21564 48596 21616
rect 48648 21604 48654 21616
rect 48685 21607 48743 21613
rect 48685 21604 48697 21607
rect 48648 21576 48697 21604
rect 48648 21564 48654 21576
rect 48685 21573 48697 21576
rect 48731 21573 48743 21607
rect 48685 21567 48743 21573
rect 49142 21564 49148 21616
rect 49200 21564 49206 21616
rect 41049 21539 41107 21545
rect 41049 21536 41061 21539
rect 40512 21508 41061 21536
rect 41049 21505 41061 21508
rect 41095 21505 41107 21539
rect 41049 21499 41107 21505
rect 44269 21539 44327 21545
rect 44269 21505 44281 21539
rect 44315 21505 44327 21539
rect 44269 21499 44327 21505
rect 45002 21496 45008 21548
rect 45060 21536 45066 21548
rect 45097 21539 45155 21545
rect 45097 21536 45109 21539
rect 45060 21508 45109 21536
rect 45060 21496 45066 21508
rect 45097 21505 45109 21508
rect 45143 21505 45155 21539
rect 45097 21499 45155 21505
rect 47581 21539 47639 21545
rect 47581 21505 47593 21539
rect 47627 21536 47639 21539
rect 47670 21536 47676 21548
rect 47627 21508 47676 21536
rect 47627 21505 47639 21508
rect 47581 21499 47639 21505
rect 47670 21496 47676 21508
rect 47728 21496 47734 21548
rect 47762 21496 47768 21548
rect 47820 21536 47826 21548
rect 47857 21539 47915 21545
rect 47857 21536 47869 21539
rect 47820 21508 47869 21536
rect 47820 21496 47826 21508
rect 47857 21505 47869 21508
rect 47903 21505 47915 21539
rect 47857 21499 47915 21505
rect 47949 21539 48007 21545
rect 47949 21505 47961 21539
rect 47995 21505 48007 21539
rect 48406 21536 48412 21548
rect 48367 21508 48412 21536
rect 47949 21499 48007 21505
rect 30524 21440 33548 21468
rect 35713 21471 35771 21477
rect 30524 21428 30530 21440
rect 35713 21437 35725 21471
rect 35759 21468 35771 21471
rect 36814 21468 36820 21480
rect 35759 21440 36820 21468
rect 35759 21437 35771 21440
rect 35713 21431 35771 21437
rect 36814 21428 36820 21440
rect 36872 21428 36878 21480
rect 39298 21428 39304 21480
rect 39356 21468 39362 21480
rect 40957 21471 41015 21477
rect 40957 21468 40969 21471
rect 39356 21440 40969 21468
rect 39356 21428 39362 21440
rect 40957 21437 40969 21440
rect 41003 21437 41015 21471
rect 42610 21468 42616 21480
rect 42571 21440 42616 21468
rect 40957 21431 41015 21437
rect 42610 21428 42616 21440
rect 42668 21428 42674 21480
rect 42702 21428 42708 21480
rect 42760 21468 42766 21480
rect 44085 21471 44143 21477
rect 44085 21468 44097 21471
rect 42760 21440 44097 21468
rect 42760 21428 42766 21440
rect 44085 21437 44097 21440
rect 44131 21437 44143 21471
rect 44085 21431 44143 21437
rect 44729 21471 44787 21477
rect 44729 21437 44741 21471
rect 44775 21437 44787 21471
rect 44729 21431 44787 21437
rect 27249 21403 27307 21409
rect 27249 21369 27261 21403
rect 27295 21369 27307 21403
rect 27249 21363 27307 21369
rect 27338 21360 27344 21412
rect 27396 21400 27402 21412
rect 27396 21372 27441 21400
rect 27396 21360 27402 21372
rect 27522 21360 27528 21412
rect 27580 21400 27586 21412
rect 29362 21400 29368 21412
rect 27580 21372 29368 21400
rect 27580 21360 27586 21372
rect 29362 21360 29368 21372
rect 29420 21360 29426 21412
rect 31846 21400 31852 21412
rect 29564 21372 31852 21400
rect 21266 21332 21272 21344
rect 19352 21304 21272 21332
rect 21266 21292 21272 21304
rect 21324 21332 21330 21344
rect 21634 21332 21640 21344
rect 21324 21304 21640 21332
rect 21324 21292 21330 21304
rect 21634 21292 21640 21304
rect 21692 21292 21698 21344
rect 22373 21335 22431 21341
rect 22373 21301 22385 21335
rect 22419 21332 22431 21335
rect 22462 21332 22468 21344
rect 22419 21304 22468 21332
rect 22419 21301 22431 21304
rect 22373 21295 22431 21301
rect 22462 21292 22468 21304
rect 22520 21332 22526 21344
rect 24946 21332 24952 21344
rect 22520 21304 24952 21332
rect 22520 21292 22526 21304
rect 24946 21292 24952 21304
rect 25004 21292 25010 21344
rect 25041 21335 25099 21341
rect 25041 21301 25053 21335
rect 25087 21332 25099 21335
rect 26234 21332 26240 21344
rect 25087 21304 26240 21332
rect 25087 21301 25099 21304
rect 25041 21295 25099 21301
rect 26234 21292 26240 21304
rect 26292 21292 26298 21344
rect 26421 21335 26479 21341
rect 26421 21301 26433 21335
rect 26467 21332 26479 21335
rect 27614 21332 27620 21344
rect 26467 21304 27620 21332
rect 26467 21301 26479 21304
rect 26421 21295 26479 21301
rect 27614 21292 27620 21304
rect 27672 21292 27678 21344
rect 27798 21292 27804 21344
rect 27856 21332 27862 21344
rect 28810 21332 28816 21344
rect 27856 21304 28816 21332
rect 27856 21292 27862 21304
rect 28810 21292 28816 21304
rect 28868 21332 28874 21344
rect 29564 21332 29592 21372
rect 31846 21360 31852 21372
rect 31904 21360 31910 21412
rect 41417 21403 41475 21409
rect 41417 21369 41429 21403
rect 41463 21400 41475 21403
rect 43622 21400 43628 21412
rect 41463 21372 43628 21400
rect 41463 21369 41475 21372
rect 41417 21363 41475 21369
rect 43622 21360 43628 21372
rect 43680 21360 43686 21412
rect 28868 21304 29592 21332
rect 28868 21292 28874 21304
rect 29822 21292 29828 21344
rect 29880 21332 29886 21344
rect 31113 21335 31171 21341
rect 31113 21332 31125 21335
rect 29880 21304 31125 21332
rect 29880 21292 29886 21304
rect 31113 21301 31125 21304
rect 31159 21301 31171 21335
rect 31113 21295 31171 21301
rect 32030 21292 32036 21344
rect 32088 21332 32094 21344
rect 32677 21335 32735 21341
rect 32677 21332 32689 21335
rect 32088 21304 32689 21332
rect 32088 21292 32094 21304
rect 32677 21301 32689 21304
rect 32723 21301 32735 21335
rect 33410 21332 33416 21344
rect 33371 21304 33416 21332
rect 32677 21295 32735 21301
rect 33410 21292 33416 21304
rect 33468 21292 33474 21344
rect 35802 21292 35808 21344
rect 35860 21332 35866 21344
rect 37369 21335 37427 21341
rect 37369 21332 37381 21335
rect 35860 21304 37381 21332
rect 35860 21292 35866 21304
rect 37369 21301 37381 21304
rect 37415 21301 37427 21335
rect 37369 21295 37427 21301
rect 43438 21292 43444 21344
rect 43496 21332 43502 21344
rect 44744 21332 44772 21431
rect 47394 21428 47400 21480
rect 47452 21428 47458 21480
rect 47412 21400 47440 21428
rect 47762 21400 47768 21412
rect 47412 21372 47768 21400
rect 47762 21360 47768 21372
rect 47820 21360 47826 21412
rect 43496 21304 44772 21332
rect 43496 21292 43502 21304
rect 47394 21292 47400 21344
rect 47452 21332 47458 21344
rect 47673 21335 47731 21341
rect 47673 21332 47685 21335
rect 47452 21304 47685 21332
rect 47452 21292 47458 21304
rect 47673 21301 47685 21304
rect 47719 21301 47731 21335
rect 47964 21332 47992 21499
rect 48406 21496 48412 21508
rect 48464 21496 48470 21548
rect 50617 21539 50675 21545
rect 50617 21505 50629 21539
rect 50663 21536 50675 21539
rect 50706 21536 50712 21548
rect 50663 21508 50712 21536
rect 50663 21505 50675 21508
rect 50617 21499 50675 21505
rect 50706 21496 50712 21508
rect 50764 21496 50770 21548
rect 53009 21539 53067 21545
rect 53009 21505 53021 21539
rect 53055 21536 53067 21539
rect 53098 21536 53104 21548
rect 53055 21508 53104 21536
rect 53055 21505 53067 21508
rect 53009 21499 53067 21505
rect 53098 21496 53104 21508
rect 53156 21496 53162 21548
rect 56686 21496 56692 21548
rect 56744 21536 56750 21548
rect 56744 21508 56810 21536
rect 56744 21496 56750 21508
rect 49326 21428 49332 21480
rect 49384 21468 49390 21480
rect 50893 21471 50951 21477
rect 50893 21468 50905 21471
rect 49384 21440 50905 21468
rect 49384 21428 49390 21440
rect 50893 21437 50905 21440
rect 50939 21437 50951 21471
rect 50893 21431 50951 21437
rect 51994 21428 52000 21480
rect 52052 21468 52058 21480
rect 54294 21468 54300 21480
rect 52052 21440 54300 21468
rect 52052 21428 52058 21440
rect 54294 21428 54300 21440
rect 54352 21468 54358 21480
rect 55122 21468 55128 21480
rect 54352 21440 55128 21468
rect 54352 21428 54358 21440
rect 55122 21428 55128 21440
rect 55180 21468 55186 21480
rect 55401 21471 55459 21477
rect 55401 21468 55413 21471
rect 55180 21440 55413 21468
rect 55180 21428 55186 21440
rect 55401 21437 55413 21440
rect 55447 21437 55459 21471
rect 55401 21431 55459 21437
rect 55677 21471 55735 21477
rect 55677 21437 55689 21471
rect 55723 21468 55735 21471
rect 55766 21468 55772 21480
rect 55723 21440 55772 21468
rect 55723 21437 55735 21440
rect 55677 21431 55735 21437
rect 55766 21428 55772 21440
rect 55824 21428 55830 21480
rect 49050 21332 49056 21344
rect 47964 21304 49056 21332
rect 47673 21295 47731 21301
rect 49050 21292 49056 21304
rect 49108 21292 49114 21344
rect 52822 21332 52828 21344
rect 52783 21304 52828 21332
rect 52822 21292 52828 21304
rect 52880 21292 52886 21344
rect 55490 21292 55496 21344
rect 55548 21332 55554 21344
rect 57149 21335 57207 21341
rect 57149 21332 57161 21335
rect 55548 21304 57161 21332
rect 55548 21292 55554 21304
rect 57149 21301 57161 21304
rect 57195 21301 57207 21335
rect 57149 21295 57207 21301
rect 1104 21242 58880 21264
rect 1104 21190 8174 21242
rect 8226 21190 8238 21242
rect 8290 21190 8302 21242
rect 8354 21190 8366 21242
rect 8418 21190 8430 21242
rect 8482 21190 22622 21242
rect 22674 21190 22686 21242
rect 22738 21190 22750 21242
rect 22802 21190 22814 21242
rect 22866 21190 22878 21242
rect 22930 21190 37070 21242
rect 37122 21190 37134 21242
rect 37186 21190 37198 21242
rect 37250 21190 37262 21242
rect 37314 21190 37326 21242
rect 37378 21190 51518 21242
rect 51570 21190 51582 21242
rect 51634 21190 51646 21242
rect 51698 21190 51710 21242
rect 51762 21190 51774 21242
rect 51826 21190 58880 21242
rect 1104 21168 58880 21190
rect 2958 21088 2964 21140
rect 3016 21128 3022 21140
rect 3602 21128 3608 21140
rect 3016 21100 3608 21128
rect 3016 21088 3022 21100
rect 3602 21088 3608 21100
rect 3660 21128 3666 21140
rect 6730 21128 6736 21140
rect 3660 21100 6736 21128
rect 3660 21088 3666 21100
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 7006 21088 7012 21140
rect 7064 21128 7070 21140
rect 7929 21131 7987 21137
rect 7929 21128 7941 21131
rect 7064 21100 7941 21128
rect 7064 21088 7070 21100
rect 7929 21097 7941 21100
rect 7975 21097 7987 21131
rect 7929 21091 7987 21097
rect 11624 21100 14780 21128
rect 5442 21020 5448 21072
rect 5500 21060 5506 21072
rect 7650 21060 7656 21072
rect 5500 21032 7656 21060
rect 5500 21020 5506 21032
rect 7650 21020 7656 21032
rect 7708 21020 7714 21072
rect 3234 20952 3240 21004
rect 3292 20952 3298 21004
rect 3970 20952 3976 21004
rect 4028 20992 4034 21004
rect 6546 20992 6552 21004
rect 4028 20964 6552 20992
rect 4028 20952 4034 20964
rect 6546 20952 6552 20964
rect 6604 20952 6610 21004
rect 10318 20952 10324 21004
rect 10376 20992 10382 21004
rect 11624 21001 11652 21100
rect 14752 21060 14780 21100
rect 16114 21088 16120 21140
rect 16172 21128 16178 21140
rect 16945 21131 17003 21137
rect 16945 21128 16957 21131
rect 16172 21100 16957 21128
rect 16172 21088 16178 21100
rect 16945 21097 16957 21100
rect 16991 21097 17003 21131
rect 19426 21128 19432 21140
rect 19387 21100 19432 21128
rect 16945 21091 17003 21097
rect 19426 21088 19432 21100
rect 19484 21088 19490 21140
rect 20530 21128 20536 21140
rect 20491 21100 20536 21128
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 22094 21128 22100 21140
rect 22055 21100 22100 21128
rect 22094 21088 22100 21100
rect 22152 21088 22158 21140
rect 23658 21128 23664 21140
rect 23619 21100 23664 21128
rect 23658 21088 23664 21100
rect 23716 21088 23722 21140
rect 24394 21128 24400 21140
rect 24355 21100 24400 21128
rect 24394 21088 24400 21100
rect 24452 21088 24458 21140
rect 24946 21128 24952 21140
rect 24859 21100 24952 21128
rect 24946 21088 24952 21100
rect 25004 21128 25010 21140
rect 27062 21128 27068 21140
rect 25004 21100 27068 21128
rect 25004 21088 25010 21100
rect 27062 21088 27068 21100
rect 27120 21088 27126 21140
rect 27246 21128 27252 21140
rect 27207 21100 27252 21128
rect 27246 21088 27252 21100
rect 27304 21088 27310 21140
rect 27982 21088 27988 21140
rect 28040 21128 28046 21140
rect 28169 21131 28227 21137
rect 28169 21128 28181 21131
rect 28040 21100 28181 21128
rect 28040 21088 28046 21100
rect 28169 21097 28181 21100
rect 28215 21097 28227 21131
rect 31294 21128 31300 21140
rect 31255 21100 31300 21128
rect 28169 21091 28227 21097
rect 31294 21088 31300 21100
rect 31352 21088 31358 21140
rect 33502 21128 33508 21140
rect 33463 21100 33508 21128
rect 33502 21088 33508 21100
rect 33560 21088 33566 21140
rect 36354 21128 36360 21140
rect 36315 21100 36360 21128
rect 36354 21088 36360 21100
rect 36412 21088 36418 21140
rect 37826 21128 37832 21140
rect 37787 21100 37832 21128
rect 37826 21088 37832 21100
rect 37884 21088 37890 21140
rect 42978 21088 42984 21140
rect 43036 21128 43042 21140
rect 46198 21128 46204 21140
rect 43036 21100 46204 21128
rect 43036 21088 43042 21100
rect 46198 21088 46204 21100
rect 46256 21088 46262 21140
rect 47210 21128 47216 21140
rect 47171 21100 47216 21128
rect 47210 21088 47216 21100
rect 47268 21088 47274 21140
rect 47486 21088 47492 21140
rect 47544 21128 47550 21140
rect 49326 21128 49332 21140
rect 47544 21100 49332 21128
rect 47544 21088 47550 21100
rect 49326 21088 49332 21100
rect 49384 21088 49390 21140
rect 50614 21128 50620 21140
rect 50575 21100 50620 21128
rect 50614 21088 50620 21100
rect 50672 21088 50678 21140
rect 55490 21128 55496 21140
rect 51276 21100 55496 21128
rect 17126 21060 17132 21072
rect 14752 21032 17132 21060
rect 17126 21020 17132 21032
rect 17184 21020 17190 21072
rect 19610 21020 19616 21072
rect 19668 21060 19674 21072
rect 19668 21032 20668 21060
rect 19668 21020 19674 21032
rect 11609 20995 11667 21001
rect 11609 20992 11621 20995
rect 10376 20964 11621 20992
rect 10376 20952 10382 20964
rect 11609 20961 11621 20964
rect 11655 20961 11667 20995
rect 11609 20955 11667 20961
rect 12526 20952 12532 21004
rect 12584 20992 12590 21004
rect 12584 20964 14136 20992
rect 12584 20952 12590 20964
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 3252 20924 3280 20952
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 1719 20896 3801 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4433 20927 4491 20933
rect 4433 20893 4445 20927
rect 4479 20924 4491 20927
rect 4982 20924 4988 20936
rect 4479 20896 4988 20924
rect 4479 20893 4491 20896
rect 4433 20887 4491 20893
rect 4982 20884 4988 20896
rect 5040 20884 5046 20936
rect 9398 20924 9404 20936
rect 9359 20896 9404 20924
rect 9398 20884 9404 20896
rect 9456 20884 9462 20936
rect 13357 20927 13415 20933
rect 13357 20893 13369 20927
rect 13403 20924 13415 20927
rect 13538 20924 13544 20936
rect 13403 20896 13544 20924
rect 13403 20893 13415 20896
rect 13357 20887 13415 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 14108 20933 14136 20964
rect 17034 20952 17040 21004
rect 17092 20992 17098 21004
rect 17957 20995 18015 21001
rect 17957 20992 17969 20995
rect 17092 20964 17969 20992
rect 17092 20952 17098 20964
rect 17957 20961 17969 20964
rect 18003 20961 18015 20995
rect 17957 20955 18015 20961
rect 20254 20952 20260 21004
rect 20312 20992 20318 21004
rect 20312 20964 20576 20992
rect 20312 20952 20318 20964
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 15194 20884 15200 20936
rect 15252 20924 15258 20936
rect 15657 20927 15715 20933
rect 15657 20924 15669 20927
rect 15252 20896 15669 20924
rect 15252 20884 15258 20896
rect 15657 20893 15669 20896
rect 15703 20893 15715 20927
rect 15657 20887 15715 20893
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 18049 20927 18107 20933
rect 18049 20924 18061 20927
rect 16540 20896 18061 20924
rect 16540 20884 16546 20896
rect 18049 20893 18061 20896
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 18690 20884 18696 20936
rect 18748 20924 18754 20936
rect 19337 20927 19395 20933
rect 19337 20924 19349 20927
rect 18748 20896 19349 20924
rect 18748 20884 18754 20896
rect 19337 20893 19349 20896
rect 19383 20893 19395 20927
rect 20346 20924 20352 20936
rect 20307 20896 20352 20924
rect 19337 20887 19395 20893
rect 20346 20884 20352 20896
rect 20404 20884 20410 20936
rect 20548 20933 20576 20964
rect 20533 20927 20591 20933
rect 20533 20893 20545 20927
rect 20579 20893 20591 20927
rect 20640 20924 20668 21032
rect 21082 21020 21088 21072
rect 21140 21060 21146 21072
rect 21542 21060 21548 21072
rect 21140 21032 21404 21060
rect 21503 21032 21548 21060
rect 21140 21020 21146 21032
rect 21266 20992 21272 21004
rect 21227 20964 21272 20992
rect 21266 20952 21272 20964
rect 21324 20952 21330 21004
rect 21376 20992 21404 21032
rect 21542 21020 21548 21032
rect 21600 21020 21606 21072
rect 21818 21020 21824 21072
rect 21876 21060 21882 21072
rect 22741 21063 22799 21069
rect 22741 21060 22753 21063
rect 21876 21032 22753 21060
rect 21876 21020 21882 21032
rect 22741 21029 22753 21032
rect 22787 21029 22799 21063
rect 22741 21023 22799 21029
rect 23842 21020 23848 21072
rect 23900 21060 23906 21072
rect 23900 21032 24900 21060
rect 23900 21020 23906 21032
rect 21376 20964 24808 20992
rect 21177 20927 21235 20933
rect 21177 20924 21189 20927
rect 20640 20896 21189 20924
rect 20533 20887 20591 20893
rect 21177 20893 21189 20896
rect 21223 20924 21235 20927
rect 22186 20924 22192 20936
rect 21223 20896 22192 20924
rect 21223 20893 21235 20896
rect 21177 20887 21235 20893
rect 22186 20884 22192 20896
rect 22244 20884 22250 20936
rect 22278 20884 22284 20936
rect 22336 20924 22342 20936
rect 22649 20927 22707 20933
rect 22649 20924 22661 20927
rect 22336 20896 22661 20924
rect 22336 20884 22342 20896
rect 22649 20893 22661 20896
rect 22695 20893 22707 20927
rect 23842 20924 23848 20936
rect 23803 20896 23848 20924
rect 22649 20887 22707 20893
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 24780 20933 24808 20964
rect 24872 20933 24900 21032
rect 24673 20927 24731 20933
rect 24673 20893 24685 20927
rect 24719 20893 24731 20927
rect 24673 20887 24731 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 24857 20927 24915 20933
rect 24857 20893 24869 20927
rect 24903 20893 24915 20927
rect 24857 20887 24915 20893
rect 3237 20859 3295 20865
rect 3237 20825 3249 20859
rect 3283 20856 3295 20859
rect 6641 20859 6699 20865
rect 3283 20828 4384 20856
rect 3283 20825 3295 20828
rect 3237 20819 3295 20825
rect 3881 20791 3939 20797
rect 3881 20757 3893 20791
rect 3927 20788 3939 20791
rect 4246 20788 4252 20800
rect 3927 20760 4252 20788
rect 3927 20757 3939 20760
rect 3881 20751 3939 20757
rect 4246 20748 4252 20760
rect 4304 20748 4310 20800
rect 4356 20788 4384 20828
rect 6641 20825 6653 20859
rect 6687 20825 6699 20859
rect 13081 20859 13139 20865
rect 12650 20828 13032 20856
rect 6641 20819 6699 20825
rect 5721 20791 5779 20797
rect 5721 20788 5733 20791
rect 4356 20760 5733 20788
rect 5721 20757 5733 20760
rect 5767 20788 5779 20791
rect 6656 20788 6684 20819
rect 5767 20760 6684 20788
rect 10689 20791 10747 20797
rect 5767 20757 5779 20760
rect 5721 20751 5779 20757
rect 10689 20757 10701 20791
rect 10735 20788 10747 20791
rect 10778 20788 10784 20800
rect 10735 20760 10784 20788
rect 10735 20757 10747 20760
rect 10689 20751 10747 20757
rect 10778 20748 10784 20760
rect 10836 20748 10842 20800
rect 13004 20788 13032 20828
rect 13081 20825 13093 20859
rect 13127 20856 13139 20859
rect 14642 20856 14648 20868
rect 13127 20828 14648 20856
rect 13127 20825 13139 20828
rect 13081 20819 13139 20825
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 24688 20856 24716 20887
rect 24964 20856 24992 21088
rect 26142 21020 26148 21072
rect 26200 21060 26206 21072
rect 26510 21060 26516 21072
rect 26200 21032 26372 21060
rect 26471 21032 26516 21060
rect 26200 21020 26206 21032
rect 25041 20927 25099 20933
rect 25041 20893 25053 20927
rect 25087 20924 25099 20927
rect 25222 20924 25228 20936
rect 25087 20896 25228 20924
rect 25087 20893 25099 20896
rect 25041 20887 25099 20893
rect 25222 20884 25228 20896
rect 25280 20884 25286 20936
rect 25685 20927 25743 20933
rect 25685 20893 25697 20927
rect 25731 20924 25743 20927
rect 26234 20924 26240 20936
rect 25731 20896 26240 20924
rect 25731 20893 25743 20896
rect 25685 20887 25743 20893
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 26344 20933 26372 21032
rect 26510 21020 26516 21032
rect 26568 21020 26574 21072
rect 27890 21060 27896 21072
rect 27264 21032 27896 21060
rect 26329 20927 26387 20933
rect 26329 20893 26341 20927
rect 26375 20893 26387 20927
rect 26329 20887 26387 20893
rect 27264 20856 27292 21032
rect 27890 21020 27896 21032
rect 27948 21060 27954 21072
rect 28994 21060 29000 21072
rect 27948 21032 29000 21060
rect 27948 21020 27954 21032
rect 27338 20952 27344 21004
rect 27396 20992 27402 21004
rect 28460 21001 28488 21032
rect 28994 21020 29000 21032
rect 29052 21020 29058 21072
rect 33520 21060 33548 21088
rect 33520 21032 34928 21060
rect 28353 20995 28411 21001
rect 28353 20992 28365 20995
rect 27396 20964 28365 20992
rect 27396 20952 27402 20964
rect 28353 20961 28365 20964
rect 28399 20961 28411 20995
rect 28353 20955 28411 20961
rect 28445 20995 28503 21001
rect 28445 20961 28457 20995
rect 28491 20961 28503 20995
rect 28445 20955 28503 20961
rect 28629 20995 28687 21001
rect 28629 20961 28641 20995
rect 28675 20992 28687 20995
rect 29270 20992 29276 21004
rect 28675 20964 29276 20992
rect 28675 20961 28687 20964
rect 28629 20955 28687 20961
rect 29270 20952 29276 20964
rect 29328 20952 29334 21004
rect 29822 20992 29828 21004
rect 29783 20964 29828 20992
rect 29822 20952 29828 20964
rect 29880 20952 29886 21004
rect 31754 20952 31760 21004
rect 31812 20992 31818 21004
rect 32030 20992 32036 21004
rect 31812 20964 31857 20992
rect 31991 20964 32036 20992
rect 31812 20952 31818 20964
rect 32030 20952 32036 20964
rect 32088 20952 32094 21004
rect 32398 20952 32404 21004
rect 32456 20992 32462 21004
rect 34057 20995 34115 21001
rect 34057 20992 34069 20995
rect 32456 20964 34069 20992
rect 32456 20952 32462 20964
rect 34057 20961 34069 20964
rect 34103 20961 34115 20995
rect 34057 20955 34115 20961
rect 27430 20924 27436 20936
rect 27391 20896 27436 20924
rect 27430 20884 27436 20896
rect 27488 20884 27494 20936
rect 27709 20927 27767 20933
rect 27709 20893 27721 20927
rect 27755 20893 27767 20927
rect 27709 20887 27767 20893
rect 28537 20927 28595 20933
rect 28537 20893 28549 20927
rect 28583 20924 28595 20927
rect 28718 20924 28724 20936
rect 28583 20896 28724 20924
rect 28583 20893 28595 20896
rect 28537 20887 28595 20893
rect 24688 20828 24992 20856
rect 25056 20828 27292 20856
rect 27724 20856 27752 20887
rect 28718 20884 28724 20896
rect 28776 20884 28782 20936
rect 29549 20927 29607 20933
rect 29549 20893 29561 20927
rect 29595 20893 29607 20927
rect 29549 20887 29607 20893
rect 34149 20927 34207 20933
rect 34149 20893 34161 20927
rect 34195 20924 34207 20927
rect 34606 20924 34612 20936
rect 34195 20896 34612 20924
rect 34195 20893 34207 20896
rect 34149 20887 34207 20893
rect 29564 20856 29592 20887
rect 34606 20884 34612 20896
rect 34664 20884 34670 20936
rect 34793 20927 34851 20933
rect 34793 20893 34805 20927
rect 34839 20893 34851 20927
rect 34900 20924 34928 21032
rect 35526 21020 35532 21072
rect 35584 21060 35590 21072
rect 37185 21063 37243 21069
rect 37185 21060 37197 21063
rect 35584 21032 37197 21060
rect 35584 21020 35590 21032
rect 37185 21029 37197 21032
rect 37231 21060 37243 21063
rect 40586 21060 40592 21072
rect 37231 21032 40592 21060
rect 37231 21029 37243 21032
rect 37185 21023 37243 21029
rect 40586 21020 40592 21032
rect 40644 21020 40650 21072
rect 42610 21020 42616 21072
rect 42668 21060 42674 21072
rect 43990 21060 43996 21072
rect 42668 21032 43996 21060
rect 42668 21020 42674 21032
rect 40957 20995 41015 21001
rect 40957 20961 40969 20995
rect 41003 20992 41015 20995
rect 42702 20992 42708 21004
rect 41003 20964 42708 20992
rect 41003 20961 41015 20964
rect 40957 20955 41015 20961
rect 42702 20952 42708 20964
rect 42760 20952 42766 21004
rect 43364 21001 43392 21032
rect 43990 21020 43996 21032
rect 44048 21020 44054 21072
rect 44266 21020 44272 21072
rect 44324 21060 44330 21072
rect 44818 21060 44824 21072
rect 44324 21032 44824 21060
rect 44324 21020 44330 21032
rect 44818 21020 44824 21032
rect 44876 21020 44882 21072
rect 43349 20995 43407 21001
rect 43349 20961 43361 20995
rect 43395 20961 43407 20995
rect 43622 20992 43628 21004
rect 43583 20964 43628 20992
rect 43349 20955 43407 20961
rect 43622 20952 43628 20964
rect 43680 20952 43686 21004
rect 46216 21001 46244 21088
rect 46842 21020 46848 21072
rect 46900 21060 46906 21072
rect 48225 21063 48283 21069
rect 48225 21060 48237 21063
rect 46900 21032 48237 21060
rect 46900 21020 46906 21032
rect 48225 21029 48237 21032
rect 48271 21029 48283 21063
rect 50338 21060 50344 21072
rect 48225 21023 48283 21029
rect 49344 21032 50344 21060
rect 43809 20995 43867 21001
rect 43809 20961 43821 20995
rect 43855 20992 43867 20995
rect 46201 20995 46259 21001
rect 43855 20964 45600 20992
rect 43855 20961 43867 20964
rect 43809 20955 43867 20961
rect 34977 20927 35035 20933
rect 34977 20924 34989 20927
rect 34900 20896 34989 20924
rect 34793 20887 34851 20893
rect 34977 20893 34989 20896
rect 35023 20893 35035 20927
rect 36538 20924 36544 20936
rect 36499 20896 36544 20924
rect 34977 20887 35035 20893
rect 29730 20856 29736 20868
rect 27724 20828 29736 20856
rect 14185 20791 14243 20797
rect 14185 20788 14197 20791
rect 13004 20760 14197 20788
rect 14185 20757 14197 20760
rect 14231 20757 14243 20791
rect 15194 20788 15200 20800
rect 15155 20760 15200 20788
rect 14185 20751 14243 20757
rect 15194 20748 15200 20760
rect 15252 20788 15258 20800
rect 16482 20788 16488 20800
rect 15252 20760 16488 20788
rect 15252 20748 15258 20760
rect 16482 20748 16488 20760
rect 16540 20748 16546 20800
rect 18414 20788 18420 20800
rect 18375 20760 18420 20788
rect 18414 20748 18420 20760
rect 18472 20748 18478 20800
rect 20438 20748 20444 20800
rect 20496 20788 20502 20800
rect 25056 20788 25084 20828
rect 29730 20816 29736 20828
rect 29788 20816 29794 20868
rect 30558 20816 30564 20868
rect 30616 20816 30622 20868
rect 33410 20856 33416 20868
rect 33258 20828 33416 20856
rect 33410 20816 33416 20828
rect 33468 20816 33474 20868
rect 25682 20788 25688 20800
rect 20496 20760 25084 20788
rect 25643 20760 25688 20788
rect 20496 20748 20502 20760
rect 25682 20748 25688 20760
rect 25740 20748 25746 20800
rect 27617 20791 27675 20797
rect 27617 20757 27629 20791
rect 27663 20788 27675 20791
rect 29086 20788 29092 20800
rect 27663 20760 29092 20788
rect 27663 20757 27675 20760
rect 27617 20751 27675 20757
rect 29086 20748 29092 20760
rect 29144 20748 29150 20800
rect 32858 20748 32864 20800
rect 32916 20788 32922 20800
rect 34808 20788 34836 20887
rect 36538 20884 36544 20896
rect 36596 20884 36602 20936
rect 36998 20884 37004 20936
rect 37056 20924 37062 20936
rect 37056 20896 37101 20924
rect 37056 20884 37062 20896
rect 37918 20884 37924 20936
rect 37976 20924 37982 20936
rect 38013 20927 38071 20933
rect 38013 20924 38025 20927
rect 37976 20896 38025 20924
rect 37976 20884 37982 20896
rect 38013 20893 38025 20896
rect 38059 20893 38071 20927
rect 38013 20887 38071 20893
rect 39301 20927 39359 20933
rect 39301 20893 39313 20927
rect 39347 20924 39359 20927
rect 39942 20924 39948 20936
rect 39347 20896 39948 20924
rect 39347 20893 39359 20896
rect 39301 20887 39359 20893
rect 39942 20884 39948 20896
rect 40000 20884 40006 20936
rect 40034 20884 40040 20936
rect 40092 20924 40098 20936
rect 40129 20927 40187 20933
rect 40129 20924 40141 20927
rect 40092 20896 40141 20924
rect 40092 20884 40098 20896
rect 40129 20893 40141 20896
rect 40175 20893 40187 20927
rect 40129 20887 40187 20893
rect 44174 20884 44180 20936
rect 44232 20924 44238 20936
rect 44269 20927 44327 20933
rect 44269 20924 44281 20927
rect 44232 20896 44281 20924
rect 44232 20884 44238 20896
rect 44269 20893 44281 20896
rect 44315 20893 44327 20927
rect 45281 20927 45339 20933
rect 45281 20924 45293 20927
rect 44269 20887 44327 20893
rect 44376 20896 45293 20924
rect 35805 20859 35863 20865
rect 35805 20825 35817 20859
rect 35851 20856 35863 20859
rect 35851 20828 41920 20856
rect 35851 20825 35863 20828
rect 35805 20819 35863 20825
rect 32916 20760 34836 20788
rect 32916 20748 32922 20760
rect 36538 20748 36544 20800
rect 36596 20788 36602 20800
rect 37918 20788 37924 20800
rect 36596 20760 37924 20788
rect 36596 20748 36602 20760
rect 37918 20748 37924 20760
rect 37976 20788 37982 20800
rect 38470 20788 38476 20800
rect 37976 20760 38476 20788
rect 37976 20748 37982 20760
rect 38470 20748 38476 20760
rect 38528 20748 38534 20800
rect 39117 20791 39175 20797
rect 39117 20757 39129 20791
rect 39163 20788 39175 20791
rect 41322 20788 41328 20800
rect 39163 20760 41328 20788
rect 39163 20757 39175 20760
rect 39117 20751 39175 20757
rect 41322 20748 41328 20760
rect 41380 20748 41386 20800
rect 41892 20788 41920 20828
rect 42426 20816 42432 20868
rect 42484 20856 42490 20868
rect 44082 20856 44088 20868
rect 42484 20828 44088 20856
rect 42484 20816 42490 20828
rect 44082 20816 44088 20828
rect 44140 20856 44146 20868
rect 44376 20856 44404 20896
rect 45281 20893 45293 20896
rect 45327 20893 45339 20927
rect 45281 20887 45339 20893
rect 44140 20828 44404 20856
rect 44140 20816 44146 20828
rect 44726 20816 44732 20868
rect 44784 20856 44790 20868
rect 44910 20856 44916 20868
rect 44784 20828 44916 20856
rect 44784 20816 44790 20828
rect 44910 20816 44916 20828
rect 44968 20856 44974 20868
rect 45005 20859 45063 20865
rect 45005 20856 45017 20859
rect 44968 20828 45017 20856
rect 44968 20816 44974 20828
rect 45005 20825 45017 20828
rect 45051 20825 45063 20859
rect 45572 20856 45600 20964
rect 46201 20961 46213 20995
rect 46247 20961 46259 20995
rect 49234 20992 49240 21004
rect 46201 20955 46259 20961
rect 47504 20964 49240 20992
rect 45738 20884 45744 20936
rect 45796 20924 45802 20936
rect 45925 20927 45983 20933
rect 45925 20924 45937 20927
rect 45796 20896 45937 20924
rect 45796 20884 45802 20896
rect 45925 20893 45937 20896
rect 45971 20893 45983 20927
rect 47394 20924 47400 20936
rect 47355 20896 47400 20924
rect 45925 20887 45983 20893
rect 47394 20884 47400 20896
rect 47452 20884 47458 20936
rect 47504 20933 47532 20964
rect 47489 20927 47547 20933
rect 47489 20893 47501 20927
rect 47535 20893 47547 20927
rect 47670 20924 47676 20936
rect 47631 20896 47676 20924
rect 47489 20887 47547 20893
rect 47670 20884 47676 20896
rect 47728 20884 47734 20936
rect 47762 20884 47768 20936
rect 47820 20924 47826 20936
rect 48406 20924 48412 20936
rect 47820 20896 47865 20924
rect 48367 20896 48412 20924
rect 47820 20884 47826 20896
rect 48406 20884 48412 20896
rect 48464 20884 48470 20936
rect 48608 20933 48636 20964
rect 49234 20952 49240 20964
rect 49292 20952 49298 21004
rect 48593 20927 48651 20933
rect 48593 20893 48605 20927
rect 48639 20893 48651 20927
rect 48593 20887 48651 20893
rect 48685 20927 48743 20933
rect 48685 20893 48697 20927
rect 48731 20893 48743 20927
rect 49344 20924 49372 21032
rect 50338 21020 50344 21032
rect 50396 21020 50402 21072
rect 48685 20887 48743 20893
rect 48792 20896 49372 20924
rect 49436 20964 51212 20992
rect 47412 20856 47440 20884
rect 48700 20856 48728 20887
rect 45572 20828 47348 20856
rect 47412 20828 48728 20856
rect 45005 20819 45063 20825
rect 44266 20788 44272 20800
rect 41892 20760 44272 20788
rect 44266 20748 44272 20760
rect 44324 20748 44330 20800
rect 44453 20791 44511 20797
rect 44453 20757 44465 20791
rect 44499 20788 44511 20791
rect 44634 20788 44640 20800
rect 44499 20760 44640 20788
rect 44499 20757 44511 20760
rect 44453 20751 44511 20757
rect 44634 20748 44640 20760
rect 44692 20748 44698 20800
rect 46474 20748 46480 20800
rect 46532 20788 46538 20800
rect 46661 20791 46719 20797
rect 46661 20788 46673 20791
rect 46532 20760 46673 20788
rect 46532 20748 46538 20760
rect 46661 20757 46673 20760
rect 46707 20757 46719 20791
rect 47320 20788 47348 20828
rect 48792 20788 48820 20896
rect 49050 20816 49056 20868
rect 49108 20856 49114 20868
rect 49297 20859 49355 20865
rect 49297 20856 49309 20859
rect 49108 20828 49309 20856
rect 49108 20816 49114 20828
rect 49297 20825 49309 20828
rect 49343 20856 49355 20859
rect 49436 20856 49464 20964
rect 50154 20924 50160 20936
rect 50115 20896 50160 20924
rect 50154 20884 50160 20896
rect 50212 20884 50218 20936
rect 50430 20924 50436 20936
rect 50391 20896 50436 20924
rect 50430 20884 50436 20896
rect 50488 20884 50494 20936
rect 51077 20927 51135 20933
rect 51077 20893 51089 20927
rect 51123 20924 51135 20927
rect 51184 20924 51212 20964
rect 51276 20936 51304 21100
rect 55490 21088 55496 21100
rect 55548 21088 55554 21140
rect 55766 21128 55772 21140
rect 55727 21100 55772 21128
rect 55766 21088 55772 21100
rect 55824 21088 55830 21140
rect 54205 21063 54263 21069
rect 54205 21029 54217 21063
rect 54251 21060 54263 21063
rect 54251 21032 55444 21060
rect 54251 21029 54263 21032
rect 54205 21023 54263 21029
rect 51721 20995 51779 21001
rect 51721 20961 51733 20995
rect 51767 20992 51779 20995
rect 51994 20992 52000 21004
rect 51767 20964 52000 20992
rect 51767 20961 51779 20964
rect 51721 20955 51779 20961
rect 51994 20952 52000 20964
rect 52052 20952 52058 21004
rect 52362 20952 52368 21004
rect 52420 20992 52426 21004
rect 52420 20964 53236 20992
rect 52420 20952 52426 20964
rect 51123 20896 51212 20924
rect 51123 20893 51135 20896
rect 51077 20887 51135 20893
rect 49343 20828 49464 20856
rect 49343 20825 49355 20828
rect 49297 20819 49355 20825
rect 49510 20816 49516 20868
rect 49568 20856 49574 20868
rect 50062 20856 50068 20868
rect 49568 20828 50068 20856
rect 49568 20816 49574 20828
rect 50062 20816 50068 20828
rect 50120 20816 50126 20868
rect 50249 20859 50307 20865
rect 50249 20825 50261 20859
rect 50295 20856 50307 20859
rect 51184 20856 51212 20896
rect 51258 20884 51264 20936
rect 51316 20924 51322 20936
rect 51316 20896 51409 20924
rect 51316 20884 51322 20896
rect 51994 20856 52000 20868
rect 50295 20828 51074 20856
rect 51184 20828 51304 20856
rect 51955 20828 52000 20856
rect 50295 20825 50307 20828
rect 50249 20819 50307 20825
rect 47320 20760 48820 20788
rect 46661 20751 46719 20757
rect 48866 20748 48872 20800
rect 48924 20788 48930 20800
rect 49145 20791 49203 20797
rect 49145 20788 49157 20791
rect 48924 20760 49157 20788
rect 48924 20748 48930 20760
rect 49145 20757 49157 20760
rect 49191 20757 49203 20791
rect 51046 20788 51074 20828
rect 51169 20791 51227 20797
rect 51169 20788 51181 20791
rect 51046 20760 51181 20788
rect 49145 20751 49203 20757
rect 51169 20757 51181 20760
rect 51215 20757 51227 20791
rect 51276 20788 51304 20828
rect 51994 20816 52000 20828
rect 52052 20816 52058 20868
rect 53208 20856 53236 20964
rect 53650 20952 53656 21004
rect 53708 20992 53714 21004
rect 55416 21001 55444 21032
rect 54297 20995 54355 21001
rect 54297 20992 54309 20995
rect 53708 20964 54309 20992
rect 53708 20952 53714 20964
rect 54297 20961 54309 20964
rect 54343 20961 54355 20995
rect 54297 20955 54355 20961
rect 55401 20995 55459 21001
rect 55401 20961 55413 20995
rect 55447 20961 55459 20995
rect 55401 20955 55459 20961
rect 53282 20884 53288 20936
rect 53340 20924 53346 20936
rect 54021 20927 54079 20933
rect 54021 20924 54033 20927
rect 53340 20896 54033 20924
rect 53340 20884 53346 20896
rect 54021 20893 54033 20896
rect 54067 20893 54079 20927
rect 54021 20887 54079 20893
rect 54110 20884 54116 20936
rect 54168 20924 54174 20936
rect 55490 20924 55496 20936
rect 54168 20896 54213 20924
rect 55451 20896 55496 20924
rect 54168 20884 54174 20896
rect 55490 20884 55496 20896
rect 55548 20884 55554 20936
rect 56686 20924 56692 20936
rect 56647 20896 56692 20924
rect 56686 20884 56692 20896
rect 56744 20884 56750 20936
rect 56704 20856 56732 20884
rect 53208 20842 56732 20856
rect 53222 20828 56732 20842
rect 56873 20859 56931 20865
rect 56873 20825 56885 20859
rect 56919 20856 56931 20859
rect 57330 20856 57336 20868
rect 56919 20828 57336 20856
rect 56919 20825 56931 20828
rect 56873 20819 56931 20825
rect 57330 20816 57336 20828
rect 57388 20816 57394 20868
rect 53282 20788 53288 20800
rect 51276 20760 53288 20788
rect 51169 20751 51227 20757
rect 53282 20748 53288 20760
rect 53340 20748 53346 20800
rect 53466 20788 53472 20800
rect 53427 20760 53472 20788
rect 53466 20748 53472 20760
rect 53524 20748 53530 20800
rect 1104 20698 58880 20720
rect 1104 20646 15398 20698
rect 15450 20646 15462 20698
rect 15514 20646 15526 20698
rect 15578 20646 15590 20698
rect 15642 20646 15654 20698
rect 15706 20646 29846 20698
rect 29898 20646 29910 20698
rect 29962 20646 29974 20698
rect 30026 20646 30038 20698
rect 30090 20646 30102 20698
rect 30154 20646 44294 20698
rect 44346 20646 44358 20698
rect 44410 20646 44422 20698
rect 44474 20646 44486 20698
rect 44538 20646 44550 20698
rect 44602 20646 58880 20698
rect 1104 20624 58880 20646
rect 2958 20584 2964 20596
rect 2919 20556 2964 20584
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 3602 20584 3608 20596
rect 3563 20556 3608 20584
rect 3602 20544 3608 20556
rect 3660 20544 3666 20596
rect 4525 20587 4583 20593
rect 4525 20553 4537 20587
rect 4571 20584 4583 20587
rect 4798 20584 4804 20596
rect 4571 20556 4804 20584
rect 4571 20553 4583 20556
rect 4525 20547 4583 20553
rect 4798 20544 4804 20556
rect 4856 20544 4862 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 7098 20584 7104 20596
rect 6687 20556 7104 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 7098 20544 7104 20556
rect 7156 20544 7162 20596
rect 7285 20587 7343 20593
rect 7285 20553 7297 20587
rect 7331 20584 7343 20587
rect 7374 20584 7380 20596
rect 7331 20556 7380 20584
rect 7331 20553 7343 20556
rect 7285 20547 7343 20553
rect 7374 20544 7380 20556
rect 7432 20544 7438 20596
rect 9122 20584 9128 20596
rect 9083 20556 9128 20584
rect 9122 20544 9128 20556
rect 9180 20544 9186 20596
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11790 20584 11796 20596
rect 11011 20556 11796 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 11790 20544 11796 20556
rect 11848 20544 11854 20596
rect 14458 20584 14464 20596
rect 14419 20556 14464 20584
rect 14458 20544 14464 20556
rect 14516 20584 14522 20596
rect 15013 20587 15071 20593
rect 15013 20584 15025 20587
rect 14516 20556 15025 20584
rect 14516 20544 14522 20556
rect 15013 20553 15025 20556
rect 15059 20584 15071 20587
rect 15194 20584 15200 20596
rect 15059 20556 15200 20584
rect 15059 20553 15071 20556
rect 15013 20547 15071 20553
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 20898 20584 20904 20596
rect 19392 20556 20904 20584
rect 19392 20544 19398 20556
rect 20898 20544 20904 20556
rect 20956 20584 20962 20596
rect 21358 20584 21364 20596
rect 20956 20556 21364 20584
rect 20956 20544 20962 20556
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 23753 20587 23811 20593
rect 23753 20553 23765 20587
rect 23799 20584 23811 20587
rect 24118 20584 24124 20596
rect 23799 20556 24124 20584
rect 23799 20553 23811 20556
rect 23753 20547 23811 20553
rect 24118 20544 24124 20556
rect 24176 20544 24182 20596
rect 25516 20556 26096 20584
rect 5813 20519 5871 20525
rect 5813 20485 5825 20519
rect 5859 20516 5871 20519
rect 7834 20516 7840 20528
rect 5859 20488 7840 20516
rect 5859 20485 5871 20488
rect 5813 20479 5871 20485
rect 7834 20476 7840 20488
rect 7892 20476 7898 20528
rect 9766 20476 9772 20528
rect 9824 20516 9830 20528
rect 10229 20519 10287 20525
rect 10229 20516 10241 20519
rect 9824 20488 10241 20516
rect 9824 20476 9830 20488
rect 10229 20485 10241 20488
rect 10275 20485 10287 20519
rect 13909 20519 13967 20525
rect 13909 20516 13921 20519
rect 13018 20488 13921 20516
rect 10229 20479 10287 20485
rect 13909 20485 13921 20488
rect 13955 20485 13967 20519
rect 13909 20479 13967 20485
rect 16758 20476 16764 20528
rect 16816 20516 16822 20528
rect 16816 20488 17816 20516
rect 16816 20476 16822 20488
rect 1949 20451 2007 20457
rect 1949 20417 1961 20451
rect 1995 20448 2007 20451
rect 2130 20448 2136 20460
rect 1995 20420 2136 20448
rect 1995 20417 2007 20420
rect 1949 20411 2007 20417
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 2774 20408 2780 20460
rect 2832 20448 2838 20460
rect 2832 20420 2877 20448
rect 2832 20408 2838 20420
rect 6362 20408 6368 20460
rect 6420 20448 6426 20460
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6420 20420 6561 20448
rect 6420 20408 6426 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 7006 20408 7012 20460
rect 7064 20448 7070 20460
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 7064 20420 7205 20448
rect 7064 20408 7070 20420
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 7650 20408 7656 20460
rect 7708 20448 7714 20460
rect 10045 20451 10103 20457
rect 10045 20448 10057 20451
rect 7708 20420 10057 20448
rect 7708 20408 7714 20420
rect 10045 20417 10057 20420
rect 10091 20417 10103 20451
rect 10778 20448 10784 20460
rect 10739 20420 10784 20448
rect 10045 20411 10103 20417
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 11422 20408 11428 20460
rect 11480 20448 11486 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 11480 20420 11529 20448
rect 11480 20408 11486 20420
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 13998 20448 14004 20460
rect 13959 20420 14004 20448
rect 11517 20411 11575 20417
rect 13998 20408 14004 20420
rect 14056 20408 14062 20460
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20448 15991 20451
rect 16390 20448 16396 20460
rect 15979 20420 16396 20448
rect 15979 20417 15991 20420
rect 15933 20411 15991 20417
rect 16390 20408 16396 20420
rect 16448 20408 16454 20460
rect 16482 20408 16488 20460
rect 16540 20448 16546 20460
rect 17497 20451 17555 20457
rect 17497 20448 17509 20451
rect 16540 20420 17509 20448
rect 16540 20408 16546 20420
rect 17497 20417 17509 20420
rect 17543 20417 17555 20451
rect 17788 20448 17816 20488
rect 17862 20476 17868 20528
rect 17920 20516 17926 20528
rect 23014 20516 23020 20528
rect 17920 20488 19380 20516
rect 20838 20488 23020 20516
rect 17920 20476 17926 20488
rect 19352 20457 19380 20488
rect 23014 20476 23020 20488
rect 23072 20476 23078 20528
rect 25516 20516 25544 20556
rect 25682 20516 25688 20528
rect 25254 20488 25544 20516
rect 25643 20488 25688 20516
rect 25682 20476 25688 20488
rect 25740 20476 25746 20528
rect 26068 20516 26096 20556
rect 26142 20544 26148 20596
rect 26200 20584 26206 20596
rect 28350 20584 28356 20596
rect 26200 20556 28356 20584
rect 26200 20544 26206 20556
rect 28350 20544 28356 20556
rect 28408 20584 28414 20596
rect 28408 20556 29408 20584
rect 28408 20544 28414 20556
rect 27890 20516 27896 20528
rect 26068 20488 27896 20516
rect 27890 20476 27896 20488
rect 27948 20476 27954 20528
rect 28258 20476 28264 20528
rect 28316 20476 28322 20528
rect 18509 20451 18567 20457
rect 18509 20448 18521 20451
rect 17788 20420 18521 20448
rect 17497 20411 17555 20417
rect 18509 20417 18521 20420
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 19337 20451 19395 20457
rect 19337 20417 19349 20451
rect 19383 20417 19395 20451
rect 22186 20448 22192 20460
rect 22147 20420 22192 20448
rect 19337 20411 19395 20417
rect 22186 20408 22192 20420
rect 22244 20408 22250 20460
rect 25958 20408 25964 20460
rect 26016 20448 26022 20460
rect 27614 20448 27620 20460
rect 26016 20420 26061 20448
rect 27575 20420 27620 20448
rect 26016 20408 26022 20420
rect 27614 20408 27620 20420
rect 27672 20408 27678 20460
rect 28074 20408 28080 20460
rect 28132 20448 28138 20460
rect 29380 20457 29408 20556
rect 29454 20544 29460 20596
rect 29512 20584 29518 20596
rect 33873 20587 33931 20593
rect 29512 20556 31754 20584
rect 29512 20544 29518 20556
rect 30098 20476 30104 20528
rect 30156 20476 30162 20528
rect 28169 20451 28227 20457
rect 28169 20448 28181 20451
rect 28132 20420 28181 20448
rect 28132 20408 28138 20420
rect 28169 20417 28181 20420
rect 28215 20417 28227 20451
rect 28169 20411 28227 20417
rect 29365 20451 29423 20457
rect 29365 20417 29377 20451
rect 29411 20417 29423 20451
rect 31726 20448 31754 20556
rect 33873 20553 33885 20587
rect 33919 20584 33931 20587
rect 39761 20587 39819 20593
rect 33919 20556 37412 20584
rect 33919 20553 33931 20556
rect 33873 20547 33931 20553
rect 32398 20516 32404 20528
rect 32359 20488 32404 20516
rect 32398 20476 32404 20488
rect 32456 20476 32462 20528
rect 32950 20476 32956 20528
rect 33008 20476 33014 20528
rect 35802 20476 35808 20528
rect 35860 20476 35866 20528
rect 36449 20519 36507 20525
rect 36449 20485 36461 20519
rect 36495 20516 36507 20519
rect 37277 20519 37335 20525
rect 37277 20516 37289 20519
rect 36495 20488 37289 20516
rect 36495 20485 36507 20488
rect 36449 20479 36507 20485
rect 37277 20485 37289 20488
rect 37323 20485 37335 20519
rect 37277 20479 37335 20485
rect 32125 20451 32183 20457
rect 32125 20448 32137 20451
rect 31726 20420 32137 20448
rect 29365 20411 29423 20417
rect 32125 20417 32137 20420
rect 32171 20417 32183 20451
rect 34514 20448 34520 20460
rect 34475 20420 34520 20448
rect 32125 20411 32183 20417
rect 34514 20408 34520 20420
rect 34572 20408 34578 20460
rect 37384 20457 37412 20556
rect 39761 20553 39773 20587
rect 39807 20584 39819 20587
rect 39942 20584 39948 20596
rect 39807 20556 39948 20584
rect 39807 20553 39819 20556
rect 39761 20547 39819 20553
rect 39942 20544 39948 20556
rect 40000 20544 40006 20596
rect 49970 20584 49976 20596
rect 48056 20556 49976 20584
rect 38746 20476 38752 20528
rect 38804 20476 38810 20528
rect 43346 20516 43352 20528
rect 42444 20488 43352 20516
rect 37369 20451 37427 20457
rect 37369 20417 37381 20451
rect 37415 20448 37427 20451
rect 37458 20448 37464 20460
rect 37415 20420 37464 20448
rect 37415 20417 37427 20420
rect 37369 20411 37427 20417
rect 37458 20408 37464 20420
rect 37516 20408 37522 20460
rect 40310 20448 40316 20460
rect 40271 20420 40316 20448
rect 40310 20408 40316 20420
rect 40368 20408 40374 20460
rect 40586 20408 40592 20460
rect 40644 20448 40650 20460
rect 42444 20457 42472 20488
rect 43346 20476 43352 20488
rect 43404 20476 43410 20528
rect 41141 20451 41199 20457
rect 41141 20448 41153 20451
rect 40644 20420 41153 20448
rect 40644 20408 40650 20420
rect 41141 20417 41153 20420
rect 41187 20417 41199 20451
rect 41141 20411 41199 20417
rect 42429 20451 42487 20457
rect 42429 20417 42441 20451
rect 42475 20417 42487 20451
rect 42429 20411 42487 20417
rect 42978 20408 42984 20460
rect 43036 20448 43042 20460
rect 43073 20451 43131 20457
rect 43073 20448 43085 20451
rect 43036 20420 43085 20448
rect 43036 20408 43042 20420
rect 43073 20417 43085 20420
rect 43119 20417 43131 20451
rect 43990 20448 43996 20460
rect 43951 20420 43996 20448
rect 43073 20411 43131 20417
rect 43990 20408 43996 20420
rect 44048 20408 44054 20460
rect 44634 20448 44640 20460
rect 44595 20420 44640 20448
rect 44634 20408 44640 20420
rect 44692 20408 44698 20460
rect 45649 20451 45707 20457
rect 45649 20417 45661 20451
rect 45695 20448 45707 20451
rect 45738 20448 45744 20460
rect 45695 20420 45744 20448
rect 45695 20417 45707 20420
rect 45649 20411 45707 20417
rect 45738 20408 45744 20420
rect 45796 20408 45802 20460
rect 46290 20448 46296 20460
rect 46251 20420 46296 20448
rect 46290 20408 46296 20420
rect 46348 20408 46354 20460
rect 47486 20408 47492 20460
rect 47544 20448 47550 20460
rect 47762 20448 47768 20460
rect 47544 20420 47768 20448
rect 47544 20408 47550 20420
rect 47762 20408 47768 20420
rect 47820 20448 47826 20460
rect 48056 20457 48084 20556
rect 49970 20544 49976 20556
rect 50028 20544 50034 20596
rect 50338 20544 50344 20596
rect 50396 20584 50402 20596
rect 51813 20587 51871 20593
rect 50396 20556 51074 20584
rect 50396 20544 50402 20556
rect 49602 20476 49608 20528
rect 49660 20476 49666 20528
rect 51046 20516 51074 20556
rect 51813 20553 51825 20587
rect 51859 20584 51871 20587
rect 51994 20584 52000 20596
rect 51859 20556 52000 20584
rect 51859 20553 51871 20556
rect 51813 20547 51871 20553
rect 51994 20544 52000 20556
rect 52052 20544 52058 20596
rect 52822 20544 52828 20596
rect 52880 20584 52886 20596
rect 52917 20587 52975 20593
rect 52917 20584 52929 20587
rect 52880 20556 52929 20584
rect 52880 20544 52886 20556
rect 52917 20553 52929 20556
rect 52963 20553 52975 20587
rect 53282 20584 53288 20596
rect 53243 20556 53288 20584
rect 52917 20547 52975 20553
rect 53282 20544 53288 20556
rect 53340 20544 53346 20596
rect 54110 20544 54116 20596
rect 54168 20584 54174 20596
rect 54205 20587 54263 20593
rect 54205 20584 54217 20587
rect 54168 20556 54217 20584
rect 54168 20544 54174 20556
rect 54205 20553 54217 20556
rect 54251 20553 54263 20587
rect 54205 20547 54263 20553
rect 53009 20519 53067 20525
rect 53009 20516 53021 20519
rect 51046 20488 53021 20516
rect 51460 20457 51488 20488
rect 53009 20485 53021 20488
rect 53055 20516 53067 20519
rect 53466 20516 53472 20528
rect 53055 20488 53472 20516
rect 53055 20485 53067 20488
rect 53009 20479 53067 20485
rect 53466 20476 53472 20488
rect 53524 20516 53530 20528
rect 53745 20519 53803 20525
rect 53745 20516 53757 20519
rect 53524 20488 53757 20516
rect 53524 20476 53530 20488
rect 53745 20485 53757 20488
rect 53791 20485 53803 20519
rect 53745 20479 53803 20485
rect 48041 20451 48099 20457
rect 48041 20448 48053 20451
rect 47820 20420 48053 20448
rect 47820 20408 47826 20420
rect 48041 20417 48053 20420
rect 48087 20417 48099 20451
rect 48041 20411 48099 20417
rect 51445 20451 51503 20457
rect 51445 20417 51457 20451
rect 51491 20417 51503 20451
rect 51445 20411 51503 20417
rect 52454 20408 52460 20460
rect 52512 20448 52518 20460
rect 53101 20451 53159 20457
rect 53101 20448 53113 20451
rect 52512 20420 53113 20448
rect 52512 20408 52518 20420
rect 53101 20417 53113 20420
rect 53147 20417 53159 20451
rect 53101 20411 53159 20417
rect 2041 20383 2099 20389
rect 2041 20349 2053 20383
rect 2087 20380 2099 20383
rect 2866 20380 2872 20392
rect 2087 20352 2872 20380
rect 2087 20349 2099 20352
rect 2041 20343 2099 20349
rect 2866 20340 2872 20352
rect 2924 20380 2930 20392
rect 3786 20380 3792 20392
rect 2924 20352 3792 20380
rect 2924 20340 2930 20352
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 11790 20380 11796 20392
rect 11751 20352 11796 20380
rect 11790 20340 11796 20352
rect 11848 20340 11854 20392
rect 16025 20383 16083 20389
rect 16025 20349 16037 20383
rect 16071 20349 16083 20383
rect 16025 20343 16083 20349
rect 2317 20315 2375 20321
rect 2317 20281 2329 20315
rect 2363 20312 2375 20315
rect 7282 20312 7288 20324
rect 2363 20284 7288 20312
rect 2363 20281 2375 20284
rect 2317 20275 2375 20281
rect 7282 20272 7288 20284
rect 7340 20272 7346 20324
rect 13538 20312 13544 20324
rect 13108 20284 13544 20312
rect 8754 20204 8760 20256
rect 8812 20244 8818 20256
rect 13108 20244 13136 20284
rect 13538 20272 13544 20284
rect 13596 20272 13602 20324
rect 16040 20312 16068 20343
rect 17034 20340 17040 20392
rect 17092 20380 17098 20392
rect 17405 20383 17463 20389
rect 17405 20380 17417 20383
rect 17092 20352 17417 20380
rect 17092 20340 17098 20352
rect 17405 20349 17417 20352
rect 17451 20349 17463 20383
rect 17405 20343 17463 20349
rect 18322 20340 18328 20392
rect 18380 20380 18386 20392
rect 18417 20383 18475 20389
rect 18417 20380 18429 20383
rect 18380 20352 18429 20380
rect 18380 20340 18386 20352
rect 18417 20349 18429 20352
rect 18463 20349 18475 20383
rect 18417 20343 18475 20349
rect 18877 20383 18935 20389
rect 18877 20349 18889 20383
rect 18923 20380 18935 20383
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 18923 20352 19625 20380
rect 18923 20349 18935 20352
rect 18877 20343 18935 20349
rect 19613 20349 19625 20352
rect 19659 20349 19671 20383
rect 19613 20343 19671 20349
rect 21266 20340 21272 20392
rect 21324 20380 21330 20392
rect 22097 20383 22155 20389
rect 22097 20380 22109 20383
rect 21324 20352 22109 20380
rect 21324 20340 21330 20352
rect 22097 20349 22109 20352
rect 22143 20349 22155 20383
rect 22097 20343 22155 20349
rect 29641 20383 29699 20389
rect 29641 20349 29653 20383
rect 29687 20380 29699 20383
rect 31018 20380 31024 20392
rect 29687 20352 31024 20380
rect 29687 20349 29699 20352
rect 29641 20343 29699 20349
rect 31018 20340 31024 20352
rect 31076 20340 31082 20392
rect 36725 20383 36783 20389
rect 36725 20380 36737 20383
rect 31128 20352 36737 20380
rect 19150 20312 19156 20324
rect 16040 20284 19156 20312
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 31128 20312 31156 20352
rect 36725 20349 36737 20352
rect 36771 20380 36783 20383
rect 38013 20383 38071 20389
rect 38013 20380 38025 20383
rect 36771 20352 38025 20380
rect 36771 20349 36783 20352
rect 36725 20343 36783 20349
rect 38013 20349 38025 20352
rect 38059 20349 38071 20383
rect 38013 20343 38071 20349
rect 38289 20383 38347 20389
rect 38289 20349 38301 20383
rect 38335 20380 38347 20383
rect 39482 20380 39488 20392
rect 38335 20352 39488 20380
rect 38335 20349 38347 20352
rect 38289 20343 38347 20349
rect 39482 20340 39488 20352
rect 39540 20340 39546 20392
rect 43622 20340 43628 20392
rect 43680 20380 43686 20392
rect 43717 20383 43775 20389
rect 43717 20380 43729 20383
rect 43680 20352 43729 20380
rect 43680 20340 43686 20352
rect 43717 20349 43729 20352
rect 43763 20349 43775 20383
rect 45370 20380 45376 20392
rect 45331 20352 45376 20380
rect 43717 20343 43775 20349
rect 45370 20340 45376 20352
rect 45428 20340 45434 20392
rect 49694 20340 49700 20392
rect 49752 20380 49758 20392
rect 50157 20383 50215 20389
rect 50157 20380 50169 20383
rect 49752 20352 50169 20380
rect 49752 20340 49758 20352
rect 50157 20349 50169 20352
rect 50203 20349 50215 20383
rect 50157 20343 50215 20349
rect 50433 20383 50491 20389
rect 50433 20349 50445 20383
rect 50479 20380 50491 20383
rect 50522 20380 50528 20392
rect 50479 20352 50528 20380
rect 50479 20349 50491 20352
rect 50433 20343 50491 20349
rect 50522 20340 50528 20352
rect 50580 20340 50586 20392
rect 51350 20380 51356 20392
rect 51311 20352 51356 20380
rect 51350 20340 51356 20352
rect 51408 20340 51414 20392
rect 53116 20380 53144 20411
rect 53742 20380 53748 20392
rect 53116 20352 53748 20380
rect 53742 20340 53748 20352
rect 53800 20340 53806 20392
rect 30668 20284 31156 20312
rect 34425 20315 34483 20321
rect 8812 20216 13136 20244
rect 8812 20204 8818 20216
rect 13170 20204 13176 20256
rect 13228 20244 13234 20256
rect 13265 20247 13323 20253
rect 13265 20244 13277 20247
rect 13228 20216 13277 20244
rect 13228 20204 13234 20216
rect 13265 20213 13277 20216
rect 13311 20213 13323 20247
rect 15562 20244 15568 20256
rect 15523 20216 15568 20244
rect 13265 20207 13323 20213
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 16758 20244 16764 20256
rect 16719 20216 16764 20244
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 17770 20244 17776 20256
rect 17731 20216 17776 20244
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 21085 20247 21143 20253
rect 21085 20213 21097 20247
rect 21131 20244 21143 20247
rect 21266 20244 21272 20256
rect 21131 20216 21272 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 22557 20247 22615 20253
rect 22557 20213 22569 20247
rect 22603 20244 22615 20247
rect 23290 20244 23296 20256
rect 22603 20216 23296 20244
rect 22603 20213 22615 20216
rect 22557 20207 22615 20213
rect 23290 20204 23296 20216
rect 23348 20204 23354 20256
rect 23842 20204 23848 20256
rect 23900 20244 23906 20256
rect 24213 20247 24271 20253
rect 24213 20244 24225 20247
rect 23900 20216 24225 20244
rect 23900 20204 23906 20216
rect 24213 20213 24225 20216
rect 24259 20244 24271 20247
rect 25682 20244 25688 20256
rect 24259 20216 25688 20244
rect 24259 20213 24271 20216
rect 24213 20207 24271 20213
rect 25682 20204 25688 20216
rect 25740 20204 25746 20256
rect 27430 20204 27436 20256
rect 27488 20244 27494 20256
rect 30668 20244 30696 20284
rect 34425 20281 34437 20315
rect 34471 20312 34483 20315
rect 45388 20312 45416 20340
rect 34471 20284 35480 20312
rect 34471 20281 34483 20284
rect 34425 20275 34483 20281
rect 27488 20216 30696 20244
rect 31113 20247 31171 20253
rect 27488 20204 27494 20216
rect 31113 20213 31125 20247
rect 31159 20244 31171 20247
rect 34330 20244 34336 20256
rect 31159 20216 34336 20244
rect 31159 20213 31171 20216
rect 31113 20207 31171 20213
rect 34330 20204 34336 20216
rect 34388 20204 34394 20256
rect 34606 20204 34612 20256
rect 34664 20244 34670 20256
rect 34977 20247 35035 20253
rect 34977 20244 34989 20247
rect 34664 20216 34989 20244
rect 34664 20204 34670 20216
rect 34977 20213 34989 20216
rect 35023 20244 35035 20247
rect 35066 20244 35072 20256
rect 35023 20216 35072 20244
rect 35023 20213 35035 20216
rect 34977 20207 35035 20213
rect 35066 20204 35072 20216
rect 35124 20204 35130 20256
rect 35452 20244 35480 20284
rect 44284 20284 45416 20312
rect 48225 20315 48283 20321
rect 39390 20244 39396 20256
rect 35452 20216 39396 20244
rect 39390 20204 39396 20216
rect 39448 20204 39454 20256
rect 40126 20204 40132 20256
rect 40184 20244 40190 20256
rect 40313 20247 40371 20253
rect 40313 20244 40325 20247
rect 40184 20216 40325 20244
rect 40184 20204 40190 20216
rect 40313 20213 40325 20216
rect 40359 20213 40371 20247
rect 41230 20244 41236 20256
rect 41191 20216 41236 20244
rect 40313 20207 40371 20213
rect 41230 20204 41236 20216
rect 41288 20204 41294 20256
rect 41782 20244 41788 20256
rect 41743 20216 41788 20244
rect 41782 20204 41788 20216
rect 41840 20204 41846 20256
rect 42426 20204 42432 20256
rect 42484 20244 42490 20256
rect 42613 20247 42671 20253
rect 42613 20244 42625 20247
rect 42484 20216 42625 20244
rect 42484 20204 42490 20216
rect 42613 20213 42625 20216
rect 42659 20213 42671 20247
rect 42613 20207 42671 20213
rect 43070 20204 43076 20256
rect 43128 20244 43134 20256
rect 43257 20247 43315 20253
rect 43257 20244 43269 20247
rect 43128 20216 43269 20244
rect 43128 20204 43134 20216
rect 43257 20213 43269 20216
rect 43303 20244 43315 20247
rect 44284 20244 44312 20284
rect 48225 20281 48237 20315
rect 48271 20312 48283 20315
rect 48406 20312 48412 20324
rect 48271 20284 48412 20312
rect 48271 20281 48283 20284
rect 48225 20275 48283 20281
rect 48406 20272 48412 20284
rect 48464 20312 48470 20324
rect 48464 20284 48820 20312
rect 48464 20272 48470 20284
rect 43303 20216 44312 20244
rect 43303 20213 43315 20216
rect 43257 20207 43315 20213
rect 44726 20204 44732 20256
rect 44784 20244 44790 20256
rect 44821 20247 44879 20253
rect 44821 20244 44833 20247
rect 44784 20216 44833 20244
rect 44784 20204 44790 20216
rect 44821 20213 44833 20216
rect 44867 20213 44879 20247
rect 44821 20207 44879 20213
rect 46477 20247 46535 20253
rect 46477 20213 46489 20247
rect 46523 20244 46535 20247
rect 46566 20244 46572 20256
rect 46523 20216 46572 20244
rect 46523 20213 46535 20216
rect 46477 20207 46535 20213
rect 46566 20204 46572 20216
rect 46624 20204 46630 20256
rect 48682 20244 48688 20256
rect 48643 20216 48688 20244
rect 48682 20204 48688 20216
rect 48740 20204 48746 20256
rect 48792 20244 48820 20284
rect 52086 20272 52092 20324
rect 52144 20312 52150 20324
rect 52733 20315 52791 20321
rect 52733 20312 52745 20315
rect 52144 20284 52745 20312
rect 52144 20272 52150 20284
rect 52733 20281 52745 20284
rect 52779 20281 52791 20315
rect 52733 20275 52791 20281
rect 53834 20272 53840 20324
rect 53892 20312 53898 20324
rect 54021 20315 54079 20321
rect 54021 20312 54033 20315
rect 53892 20284 54033 20312
rect 53892 20272 53898 20284
rect 54021 20281 54033 20284
rect 54067 20281 54079 20315
rect 54021 20275 54079 20281
rect 50430 20244 50436 20256
rect 48792 20216 50436 20244
rect 50430 20204 50436 20216
rect 50488 20244 50494 20256
rect 52914 20244 52920 20256
rect 50488 20216 52920 20244
rect 50488 20204 50494 20216
rect 52914 20204 52920 20216
rect 52972 20244 52978 20256
rect 55214 20244 55220 20256
rect 52972 20216 55220 20244
rect 52972 20204 52978 20216
rect 55214 20204 55220 20216
rect 55272 20204 55278 20256
rect 1104 20154 58880 20176
rect 1104 20102 8174 20154
rect 8226 20102 8238 20154
rect 8290 20102 8302 20154
rect 8354 20102 8366 20154
rect 8418 20102 8430 20154
rect 8482 20102 22622 20154
rect 22674 20102 22686 20154
rect 22738 20102 22750 20154
rect 22802 20102 22814 20154
rect 22866 20102 22878 20154
rect 22930 20102 37070 20154
rect 37122 20102 37134 20154
rect 37186 20102 37198 20154
rect 37250 20102 37262 20154
rect 37314 20102 37326 20154
rect 37378 20102 51518 20154
rect 51570 20102 51582 20154
rect 51634 20102 51646 20154
rect 51698 20102 51710 20154
rect 51762 20102 51774 20154
rect 51826 20102 58880 20154
rect 1104 20080 58880 20102
rect 3053 20043 3111 20049
rect 3053 20009 3065 20043
rect 3099 20040 3111 20043
rect 7926 20040 7932 20052
rect 3099 20012 7932 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 10410 20040 10416 20052
rect 10183 20012 10416 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 10410 20000 10416 20012
rect 10468 20000 10474 20052
rect 10781 20043 10839 20049
rect 10781 20009 10793 20043
rect 10827 20040 10839 20043
rect 13906 20040 13912 20052
rect 10827 20012 13912 20040
rect 10827 20009 10839 20012
rect 10781 20003 10839 20009
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 18601 20043 18659 20049
rect 18601 20040 18613 20043
rect 17920 20012 18613 20040
rect 17920 20000 17926 20012
rect 18601 20009 18613 20012
rect 18647 20009 18659 20043
rect 18601 20003 18659 20009
rect 20898 20000 20904 20052
rect 20956 20040 20962 20052
rect 20956 20012 22324 20040
rect 20956 20000 20962 20012
rect 2501 19975 2559 19981
rect 2501 19941 2513 19975
rect 2547 19972 2559 19975
rect 3878 19972 3884 19984
rect 2547 19944 3884 19972
rect 2547 19941 2559 19944
rect 2501 19935 2559 19941
rect 3878 19932 3884 19944
rect 3936 19932 3942 19984
rect 5718 19932 5724 19984
rect 5776 19972 5782 19984
rect 6457 19975 6515 19981
rect 6457 19972 6469 19975
rect 5776 19944 6469 19972
rect 5776 19932 5782 19944
rect 6457 19941 6469 19944
rect 6503 19941 6515 19975
rect 15562 19972 15568 19984
rect 6457 19935 6515 19941
rect 9416 19944 11376 19972
rect 2222 19904 2228 19916
rect 2183 19876 2228 19904
rect 2222 19864 2228 19876
rect 2280 19864 2286 19916
rect 9122 19904 9128 19916
rect 5920 19876 9128 19904
rect 2130 19836 2136 19848
rect 2091 19808 2136 19836
rect 2130 19796 2136 19808
rect 2188 19796 2194 19848
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3694 19836 3700 19848
rect 3191 19808 3700 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 5920 19845 5948 19876
rect 9122 19864 9128 19876
rect 9180 19864 9186 19916
rect 5905 19839 5963 19845
rect 5905 19805 5917 19839
rect 5951 19805 5963 19839
rect 5905 19799 5963 19805
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 9416 19836 9444 19944
rect 11238 19904 11244 19916
rect 11199 19876 11244 19904
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 11348 19904 11376 19944
rect 12544 19944 15568 19972
rect 12544 19904 12572 19944
rect 15562 19932 15568 19944
rect 15620 19932 15626 19984
rect 18322 19932 18328 19984
rect 18380 19972 18386 19984
rect 20533 19975 20591 19981
rect 20533 19972 20545 19975
rect 18380 19944 20545 19972
rect 18380 19932 18386 19944
rect 20533 19941 20545 19944
rect 20579 19941 20591 19975
rect 22186 19972 22192 19984
rect 22147 19944 22192 19972
rect 20533 19935 20591 19941
rect 22186 19932 22192 19944
rect 22244 19932 22250 19984
rect 22296 19972 22324 20012
rect 22370 20000 22376 20052
rect 22428 20040 22434 20052
rect 25038 20040 25044 20052
rect 22428 20012 25044 20040
rect 22428 20000 22434 20012
rect 25038 20000 25044 20012
rect 25096 20000 25102 20052
rect 25130 20000 25136 20052
rect 25188 20040 25194 20052
rect 28905 20043 28963 20049
rect 25188 20012 26234 20040
rect 25188 20000 25194 20012
rect 26206 19972 26234 20012
rect 28905 20009 28917 20043
rect 28951 20040 28963 20043
rect 30098 20040 30104 20052
rect 28951 20012 30104 20040
rect 28951 20009 28963 20012
rect 28905 20003 28963 20009
rect 30098 20000 30104 20012
rect 30156 20000 30162 20052
rect 32950 20040 32956 20052
rect 32911 20012 32956 20040
rect 32950 20000 32956 20012
rect 33008 20000 33014 20052
rect 35452 20012 38700 20040
rect 27614 19972 27620 19984
rect 22296 19944 25636 19972
rect 26206 19944 27620 19972
rect 11348 19876 12572 19904
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 16482 19904 16488 19916
rect 12768 19876 15792 19904
rect 16443 19876 16488 19904
rect 12768 19864 12774 19876
rect 8251 19808 9444 19836
rect 9493 19839 9551 19845
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 9493 19805 9505 19839
rect 9539 19805 9551 19839
rect 9493 19799 9551 19805
rect 6270 19728 6276 19780
rect 6328 19768 6334 19780
rect 6328 19740 6762 19768
rect 6328 19728 6334 19740
rect 7650 19728 7656 19780
rect 7708 19768 7714 19780
rect 7929 19771 7987 19777
rect 7929 19768 7941 19771
rect 7708 19740 7941 19768
rect 7708 19728 7714 19740
rect 7929 19737 7941 19740
rect 7975 19737 7987 19771
rect 9508 19768 9536 19799
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9916 19808 9965 19836
rect 9916 19796 9922 19808
rect 9953 19805 9965 19808
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 10226 19796 10232 19848
rect 10284 19836 10290 19848
rect 10597 19839 10655 19845
rect 10597 19836 10609 19839
rect 10284 19808 10609 19836
rect 10284 19796 10290 19808
rect 10597 19805 10609 19808
rect 10643 19836 10655 19839
rect 10778 19836 10784 19848
rect 10643 19808 10784 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 10778 19796 10784 19808
rect 10836 19796 10842 19848
rect 14090 19796 14096 19848
rect 14148 19836 14154 19848
rect 15764 19845 15792 19876
rect 16482 19864 16488 19876
rect 16540 19864 16546 19916
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 19426 19864 19432 19876
rect 19484 19904 19490 19916
rect 20438 19904 20444 19916
rect 19484 19876 20444 19904
rect 19484 19864 19490 19876
rect 20438 19864 20444 19876
rect 20496 19904 20502 19916
rect 21545 19907 21603 19913
rect 21545 19904 21557 19907
rect 20496 19876 21557 19904
rect 20496 19864 20502 19876
rect 21545 19873 21557 19876
rect 21591 19873 21603 19907
rect 21545 19867 21603 19873
rect 22649 19907 22707 19913
rect 22649 19873 22661 19907
rect 22695 19904 22707 19907
rect 24854 19904 24860 19916
rect 22695 19876 24860 19904
rect 22695 19873 22707 19876
rect 22649 19867 22707 19873
rect 24854 19864 24860 19876
rect 24912 19864 24918 19916
rect 14829 19839 14887 19845
rect 14829 19836 14841 19839
rect 14148 19808 14841 19836
rect 14148 19796 14154 19808
rect 14829 19805 14841 19808
rect 14875 19805 14887 19839
rect 14829 19799 14887 19805
rect 15565 19839 15623 19845
rect 15565 19805 15577 19839
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19805 15807 19839
rect 17126 19836 17132 19848
rect 17087 19808 17132 19836
rect 15749 19799 15807 19805
rect 9508 19740 11008 19768
rect 7929 19731 7987 19737
rect 4617 19703 4675 19709
rect 4617 19669 4629 19703
rect 4663 19700 4675 19703
rect 5626 19700 5632 19712
rect 4663 19672 5632 19700
rect 4663 19669 4675 19672
rect 4617 19663 4675 19669
rect 5626 19660 5632 19672
rect 5684 19700 5690 19712
rect 6362 19700 6368 19712
rect 5684 19672 6368 19700
rect 5684 19660 5690 19672
rect 6362 19660 6368 19672
rect 6420 19660 6426 19712
rect 9401 19703 9459 19709
rect 9401 19669 9413 19703
rect 9447 19700 9459 19703
rect 9766 19700 9772 19712
rect 9447 19672 9772 19700
rect 9447 19669 9459 19672
rect 9401 19663 9459 19669
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 10980 19700 11008 19740
rect 11054 19728 11060 19780
rect 11112 19768 11118 19780
rect 11517 19771 11575 19777
rect 11517 19768 11529 19771
rect 11112 19740 11529 19768
rect 11112 19728 11118 19740
rect 11517 19737 11529 19740
rect 11563 19737 11575 19771
rect 11517 19731 11575 19737
rect 12526 19728 12532 19780
rect 12584 19728 12590 19780
rect 15580 19768 15608 19799
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 12912 19740 15608 19768
rect 11606 19700 11612 19712
rect 10980 19672 11612 19700
rect 11606 19660 11612 19672
rect 11664 19700 11670 19712
rect 12912 19700 12940 19740
rect 11664 19672 12940 19700
rect 12989 19703 13047 19709
rect 11664 19660 11670 19672
rect 12989 19669 13001 19703
rect 13035 19700 13047 19703
rect 13354 19700 13360 19712
rect 13035 19672 13360 19700
rect 13035 19669 13047 19672
rect 12989 19663 13047 19669
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 14366 19700 14372 19712
rect 13596 19672 14372 19700
rect 13596 19660 13602 19672
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 14550 19700 14556 19712
rect 14511 19672 14556 19700
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 14734 19660 14740 19712
rect 14792 19700 14798 19712
rect 17328 19700 17356 19799
rect 17402 19728 17408 19780
rect 17460 19768 17466 19780
rect 19536 19768 19564 19799
rect 19610 19796 19616 19848
rect 19668 19836 19674 19848
rect 20349 19839 20407 19845
rect 20349 19836 20361 19839
rect 19668 19808 20361 19836
rect 19668 19796 19674 19808
rect 20349 19805 20361 19808
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 20533 19839 20591 19845
rect 20533 19805 20545 19839
rect 20579 19836 20591 19839
rect 20898 19836 20904 19848
rect 20579 19808 20904 19836
rect 20579 19805 20591 19808
rect 20533 19799 20591 19805
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 21266 19836 21272 19848
rect 21227 19808 21272 19836
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 22462 19796 22468 19848
rect 22520 19836 22526 19848
rect 25608 19845 25636 19944
rect 27614 19932 27620 19944
rect 27672 19932 27678 19984
rect 27890 19932 27896 19984
rect 27948 19972 27954 19984
rect 29641 19975 29699 19981
rect 29641 19972 29653 19975
rect 27948 19944 29653 19972
rect 27948 19932 27954 19944
rect 29641 19941 29653 19944
rect 29687 19941 29699 19975
rect 29641 19935 29699 19941
rect 25682 19864 25688 19916
rect 25740 19904 25746 19916
rect 32401 19907 32459 19913
rect 25740 19876 26556 19904
rect 25740 19864 25746 19876
rect 22557 19839 22615 19845
rect 22557 19836 22569 19839
rect 22520 19808 22569 19836
rect 22520 19796 22526 19808
rect 22557 19805 22569 19808
rect 22603 19836 22615 19839
rect 23201 19839 23259 19845
rect 23201 19836 23213 19839
rect 22603 19808 23213 19836
rect 22603 19805 22615 19808
rect 22557 19799 22615 19805
rect 23201 19805 23213 19808
rect 23247 19805 23259 19839
rect 25593 19839 25651 19845
rect 23201 19799 23259 19805
rect 23308 19808 24900 19836
rect 20622 19768 20628 19780
rect 17460 19740 20628 19768
rect 17460 19728 17466 19740
rect 20622 19728 20628 19740
rect 20680 19728 20686 19780
rect 22278 19728 22284 19780
rect 22336 19768 22342 19780
rect 23014 19768 23020 19780
rect 22336 19740 23020 19768
rect 22336 19728 22342 19740
rect 23014 19728 23020 19740
rect 23072 19768 23078 19780
rect 23308 19768 23336 19808
rect 24872 19777 24900 19808
rect 25593 19805 25605 19839
rect 25639 19805 25651 19839
rect 25593 19799 25651 19805
rect 25777 19839 25835 19845
rect 25777 19805 25789 19839
rect 25823 19836 25835 19839
rect 25866 19836 25872 19848
rect 25823 19808 25872 19836
rect 25823 19805 25835 19808
rect 25777 19799 25835 19805
rect 25866 19796 25872 19808
rect 25924 19796 25930 19848
rect 26234 19796 26240 19848
rect 26292 19836 26298 19848
rect 26528 19845 26556 19876
rect 32401 19873 32413 19907
rect 32447 19904 32459 19907
rect 32447 19876 33732 19904
rect 32447 19873 32459 19876
rect 32401 19867 32459 19873
rect 26329 19839 26387 19845
rect 26329 19836 26341 19839
rect 26292 19808 26341 19836
rect 26292 19796 26298 19808
rect 26329 19805 26341 19808
rect 26375 19805 26387 19839
rect 26329 19799 26387 19805
rect 26513 19839 26571 19845
rect 26513 19805 26525 19839
rect 26559 19805 26571 19839
rect 26513 19799 26571 19805
rect 27890 19796 27896 19848
rect 27948 19836 27954 19848
rect 28258 19836 28264 19848
rect 27948 19808 28264 19836
rect 27948 19796 27954 19808
rect 28258 19796 28264 19808
rect 28316 19796 28322 19848
rect 28810 19836 28816 19848
rect 28771 19808 28816 19836
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 29733 19839 29791 19845
rect 29733 19805 29745 19839
rect 29779 19836 29791 19839
rect 30466 19836 30472 19848
rect 29779 19808 30472 19836
rect 29779 19805 29791 19808
rect 29733 19799 29791 19805
rect 30466 19796 30472 19808
rect 30524 19796 30530 19848
rect 30650 19836 30656 19848
rect 30611 19808 30656 19836
rect 30650 19796 30656 19808
rect 30708 19796 30714 19848
rect 33704 19845 33732 19876
rect 32861 19839 32919 19845
rect 32861 19805 32873 19839
rect 32907 19805 32919 19839
rect 32861 19799 32919 19805
rect 33689 19839 33747 19845
rect 33689 19805 33701 19839
rect 33735 19836 33747 19839
rect 34606 19836 34612 19848
rect 33735 19808 34612 19836
rect 33735 19805 33747 19808
rect 33689 19799 33747 19805
rect 23072 19740 23336 19768
rect 24857 19771 24915 19777
rect 23072 19728 23078 19740
rect 24857 19737 24869 19771
rect 24903 19737 24915 19771
rect 24857 19731 24915 19737
rect 25041 19771 25099 19777
rect 25041 19737 25053 19771
rect 25087 19768 25099 19771
rect 25130 19768 25136 19780
rect 25087 19740 25136 19768
rect 25087 19737 25099 19740
rect 25041 19731 25099 19737
rect 25130 19728 25136 19740
rect 25188 19728 25194 19780
rect 25685 19771 25743 19777
rect 25685 19737 25697 19771
rect 25731 19768 25743 19771
rect 27798 19768 27804 19780
rect 25731 19740 27660 19768
rect 27759 19740 27804 19768
rect 25731 19737 25743 19740
rect 25685 19731 25743 19737
rect 14792 19672 17356 19700
rect 18141 19703 18199 19709
rect 14792 19660 14798 19672
rect 18141 19669 18153 19703
rect 18187 19700 18199 19703
rect 19242 19700 19248 19712
rect 18187 19672 19248 19700
rect 18187 19669 18199 19672
rect 18141 19663 18199 19669
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 19886 19700 19892 19712
rect 19847 19672 19892 19700
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 23750 19700 23756 19712
rect 23711 19672 23756 19700
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 27338 19700 27344 19712
rect 27299 19672 27344 19700
rect 27338 19660 27344 19672
rect 27396 19660 27402 19712
rect 27632 19700 27660 19740
rect 27798 19728 27804 19740
rect 27856 19728 27862 19780
rect 28169 19771 28227 19777
rect 28169 19737 28181 19771
rect 28215 19768 28227 19771
rect 28994 19768 29000 19780
rect 28215 19740 29000 19768
rect 28215 19737 28227 19740
rect 28169 19731 28227 19737
rect 28994 19728 29000 19740
rect 29052 19728 29058 19780
rect 30929 19771 30987 19777
rect 30929 19737 30941 19771
rect 30975 19768 30987 19771
rect 31202 19768 31208 19780
rect 30975 19740 31208 19768
rect 30975 19737 30987 19740
rect 30929 19731 30987 19737
rect 31202 19728 31208 19740
rect 31260 19728 31266 19780
rect 31938 19728 31944 19780
rect 31996 19728 32002 19780
rect 32876 19768 32904 19799
rect 34606 19796 34612 19808
rect 34664 19796 34670 19848
rect 35452 19768 35480 20012
rect 38672 19981 38700 20012
rect 38838 20000 38844 20052
rect 38896 20040 38902 20052
rect 39853 20043 39911 20049
rect 38896 20012 39528 20040
rect 38896 20000 38902 20012
rect 38657 19975 38715 19981
rect 38657 19941 38669 19975
rect 38703 19972 38715 19975
rect 39500 19972 39528 20012
rect 39853 20009 39865 20043
rect 39899 20040 39911 20043
rect 40034 20040 40040 20052
rect 39899 20012 40040 20040
rect 39899 20009 39911 20012
rect 39853 20003 39911 20009
rect 40034 20000 40040 20012
rect 40092 20000 40098 20052
rect 40678 20040 40684 20052
rect 40144 20012 40684 20040
rect 40144 19972 40172 20012
rect 40678 20000 40684 20012
rect 40736 20040 40742 20052
rect 42610 20040 42616 20052
rect 40736 20012 42616 20040
rect 40736 20000 40742 20012
rect 42610 20000 42616 20012
rect 42668 20040 42674 20052
rect 42705 20043 42763 20049
rect 42705 20040 42717 20043
rect 42668 20012 42717 20040
rect 42668 20000 42674 20012
rect 42705 20009 42717 20012
rect 42751 20009 42763 20043
rect 43622 20040 43628 20052
rect 42705 20003 42763 20009
rect 43272 20012 43628 20040
rect 38703 19944 39436 19972
rect 39500 19944 40172 19972
rect 38703 19941 38715 19944
rect 38657 19935 38715 19941
rect 39408 19904 39436 19944
rect 41690 19932 41696 19984
rect 41748 19972 41754 19984
rect 42245 19975 42303 19981
rect 42245 19972 42257 19975
rect 41748 19944 42257 19972
rect 41748 19932 41754 19944
rect 42245 19941 42257 19944
rect 42291 19941 42303 19975
rect 42245 19935 42303 19941
rect 43272 19916 43300 20012
rect 43622 20000 43628 20012
rect 43680 20040 43686 20052
rect 50154 20040 50160 20052
rect 43680 20012 45048 20040
rect 50115 20012 50160 20040
rect 43680 20000 43686 20012
rect 40862 19904 40868 19916
rect 36648 19876 39344 19904
rect 39408 19876 40868 19904
rect 35618 19836 35624 19848
rect 35579 19808 35624 19836
rect 35618 19796 35624 19808
rect 35676 19796 35682 19848
rect 36648 19822 36676 19876
rect 38010 19796 38016 19848
rect 38068 19836 38074 19848
rect 38470 19836 38476 19848
rect 38068 19808 38113 19836
rect 38431 19808 38476 19836
rect 38068 19796 38074 19808
rect 38470 19796 38476 19808
rect 38528 19796 38534 19848
rect 37737 19771 37795 19777
rect 32416 19740 35480 19768
rect 35544 19740 36492 19768
rect 27706 19700 27712 19712
rect 27632 19672 27712 19700
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 31110 19660 31116 19712
rect 31168 19700 31174 19712
rect 32416 19700 32444 19740
rect 31168 19672 32444 19700
rect 31168 19660 31174 19672
rect 32490 19660 32496 19712
rect 32548 19700 32554 19712
rect 35544 19709 35572 19740
rect 33597 19703 33655 19709
rect 33597 19700 33609 19703
rect 32548 19672 33609 19700
rect 32548 19660 32554 19672
rect 33597 19669 33609 19672
rect 33643 19669 33655 19703
rect 33597 19663 33655 19669
rect 35529 19703 35587 19709
rect 35529 19669 35541 19703
rect 35575 19669 35587 19703
rect 36262 19700 36268 19712
rect 36223 19672 36268 19700
rect 35529 19663 35587 19669
rect 36262 19660 36268 19672
rect 36320 19660 36326 19712
rect 36464 19700 36492 19740
rect 37737 19737 37749 19771
rect 37783 19768 37795 19771
rect 38746 19768 38752 19780
rect 37783 19740 38752 19768
rect 37783 19737 37795 19740
rect 37737 19731 37795 19737
rect 38746 19728 38752 19740
rect 38804 19728 38810 19780
rect 39206 19768 39212 19780
rect 39167 19740 39212 19768
rect 39206 19728 39212 19740
rect 39264 19728 39270 19780
rect 38838 19700 38844 19712
rect 36464 19672 38844 19700
rect 38838 19660 38844 19672
rect 38896 19660 38902 19712
rect 39316 19700 39344 19876
rect 40862 19864 40868 19876
rect 40920 19864 40926 19916
rect 41322 19904 41328 19916
rect 41283 19876 41328 19904
rect 41322 19864 41328 19876
rect 41380 19864 41386 19916
rect 41601 19907 41659 19913
rect 41601 19873 41613 19907
rect 41647 19904 41659 19907
rect 41782 19904 41788 19916
rect 41647 19876 41788 19904
rect 41647 19873 41659 19876
rect 41601 19867 41659 19873
rect 41782 19864 41788 19876
rect 41840 19864 41846 19916
rect 43254 19904 43260 19916
rect 43167 19876 43260 19904
rect 43254 19864 43260 19876
rect 43312 19864 43318 19916
rect 45020 19913 45048 20012
rect 50154 20000 50160 20012
rect 50212 20000 50218 20052
rect 50338 20040 50344 20052
rect 50299 20012 50344 20040
rect 50338 20000 50344 20012
rect 50396 20000 50402 20052
rect 50430 20000 50436 20052
rect 50488 20040 50494 20052
rect 51077 20043 51135 20049
rect 51077 20040 51089 20043
rect 50488 20012 51089 20040
rect 50488 20000 50494 20012
rect 51077 20009 51089 20012
rect 51123 20009 51135 20043
rect 51077 20003 51135 20009
rect 53190 20000 53196 20052
rect 53248 20040 53254 20052
rect 53837 20043 53895 20049
rect 53837 20040 53849 20043
rect 53248 20012 53849 20040
rect 53248 20000 53254 20012
rect 53837 20009 53849 20012
rect 53883 20009 53895 20043
rect 58069 20043 58127 20049
rect 58069 20040 58081 20043
rect 53837 20003 53895 20009
rect 55600 20012 58081 20040
rect 52086 19972 52092 19984
rect 48976 19944 52092 19972
rect 48976 19913 49004 19944
rect 52086 19932 52092 19944
rect 52144 19932 52150 19984
rect 52546 19932 52552 19984
rect 52604 19972 52610 19984
rect 53650 19972 53656 19984
rect 52604 19944 53656 19972
rect 52604 19932 52610 19944
rect 53650 19932 53656 19944
rect 53708 19972 53714 19984
rect 53929 19975 53987 19981
rect 53708 19944 53880 19972
rect 53708 19932 53714 19944
rect 45005 19907 45063 19913
rect 45005 19873 45017 19907
rect 45051 19873 45063 19907
rect 45005 19867 45063 19873
rect 48961 19907 49019 19913
rect 48961 19873 48973 19907
rect 49007 19873 49019 19907
rect 50154 19904 50160 19916
rect 48961 19867 49019 19873
rect 49436 19876 50160 19904
rect 42058 19836 42064 19848
rect 42019 19808 42064 19836
rect 42058 19796 42064 19808
rect 42116 19796 42122 19848
rect 43530 19836 43536 19848
rect 43491 19808 43536 19836
rect 43530 19796 43536 19808
rect 43588 19796 43594 19848
rect 44177 19839 44235 19845
rect 44177 19805 44189 19839
rect 44223 19836 44235 19839
rect 44634 19836 44640 19848
rect 44223 19808 44640 19836
rect 44223 19805 44235 19808
rect 44177 19799 44235 19805
rect 44634 19796 44640 19808
rect 44692 19836 44698 19848
rect 45281 19839 45339 19845
rect 44692 19808 44772 19836
rect 44692 19796 44698 19808
rect 39390 19728 39396 19780
rect 39448 19768 39454 19780
rect 44453 19771 44511 19777
rect 39448 19740 40158 19768
rect 39448 19728 39454 19740
rect 44453 19737 44465 19771
rect 44499 19737 44511 19771
rect 44744 19768 44772 19808
rect 45281 19805 45293 19839
rect 45327 19836 45339 19839
rect 45738 19836 45744 19848
rect 45327 19808 45744 19836
rect 45327 19805 45339 19808
rect 45281 19799 45339 19805
rect 45738 19796 45744 19808
rect 45796 19796 45802 19848
rect 49436 19845 49464 19876
rect 50154 19864 50160 19876
rect 50212 19864 50218 19916
rect 51997 19907 52055 19913
rect 51997 19904 52009 19907
rect 50356 19876 52009 19904
rect 50356 19848 50384 19876
rect 51997 19873 52009 19876
rect 52043 19904 52055 19907
rect 52822 19904 52828 19916
rect 52043 19876 52828 19904
rect 52043 19873 52055 19876
rect 51997 19867 52055 19873
rect 52822 19864 52828 19876
rect 52880 19864 52886 19916
rect 53006 19904 53012 19916
rect 52967 19876 53012 19904
rect 53006 19864 53012 19876
rect 53064 19864 53070 19916
rect 53852 19904 53880 19944
rect 53929 19941 53941 19975
rect 53975 19972 53987 19975
rect 55600 19972 55628 20012
rect 58069 20009 58081 20012
rect 58115 20009 58127 20043
rect 58069 20003 58127 20009
rect 53975 19944 55444 19972
rect 53975 19941 53987 19944
rect 53929 19935 53987 19941
rect 55416 19913 55444 19944
rect 55508 19944 55628 19972
rect 54021 19907 54079 19913
rect 54021 19904 54033 19907
rect 53852 19876 54033 19904
rect 54021 19873 54033 19876
rect 54067 19873 54079 19907
rect 54021 19867 54079 19873
rect 55401 19907 55459 19913
rect 55401 19873 55413 19907
rect 55447 19873 55459 19907
rect 55401 19867 55459 19873
rect 45925 19839 45983 19845
rect 45925 19805 45937 19839
rect 45971 19805 45983 19839
rect 45925 19799 45983 19805
rect 49421 19839 49479 19845
rect 49421 19805 49433 19839
rect 49467 19805 49479 19839
rect 49421 19799 49479 19805
rect 49605 19839 49663 19845
rect 49605 19805 49617 19839
rect 49651 19805 49663 19839
rect 50338 19836 50344 19848
rect 50299 19808 50344 19836
rect 49605 19799 49663 19805
rect 45940 19768 45968 19799
rect 44744 19740 45968 19768
rect 46201 19771 46259 19777
rect 44453 19731 44511 19737
rect 46201 19737 46213 19771
rect 46247 19737 46259 19771
rect 46201 19731 46259 19737
rect 42150 19700 42156 19712
rect 39316 19672 42156 19700
rect 42150 19660 42156 19672
rect 42208 19660 42214 19712
rect 44468 19700 44496 19731
rect 44726 19700 44732 19712
rect 44468 19672 44732 19700
rect 44726 19660 44732 19672
rect 44784 19700 44790 19712
rect 46216 19700 46244 19731
rect 46474 19728 46480 19780
rect 46532 19768 46538 19780
rect 47121 19771 47179 19777
rect 47121 19768 47133 19771
rect 46532 19740 47133 19768
rect 46532 19728 46538 19740
rect 47121 19737 47133 19740
rect 47167 19737 47179 19771
rect 48774 19768 48780 19780
rect 48735 19740 48780 19768
rect 47121 19731 47179 19737
rect 48774 19728 48780 19740
rect 48832 19728 48838 19780
rect 49326 19728 49332 19780
rect 49384 19768 49390 19780
rect 49620 19768 49648 19799
rect 50338 19796 50344 19808
rect 50396 19796 50402 19848
rect 50430 19796 50436 19848
rect 50488 19836 50494 19848
rect 51258 19836 51264 19848
rect 50488 19808 50581 19836
rect 51219 19808 51264 19836
rect 50488 19796 50494 19808
rect 51258 19796 51264 19808
rect 51316 19796 51322 19848
rect 51905 19839 51963 19845
rect 51905 19805 51917 19839
rect 51951 19805 51963 19839
rect 52086 19836 52092 19848
rect 52048 19808 52092 19836
rect 51905 19799 51963 19805
rect 49384 19740 49648 19768
rect 49384 19728 49390 19740
rect 50062 19728 50068 19780
rect 50120 19768 50126 19780
rect 50448 19768 50476 19796
rect 50120 19740 50476 19768
rect 50617 19771 50675 19777
rect 50120 19728 50126 19740
rect 50617 19737 50629 19771
rect 50663 19768 50675 19771
rect 50798 19768 50804 19780
rect 50663 19740 50804 19768
rect 50663 19737 50675 19740
rect 50617 19731 50675 19737
rect 50798 19728 50804 19740
rect 50856 19728 50862 19780
rect 46566 19700 46572 19712
rect 44784 19672 46572 19700
rect 44784 19660 44790 19672
rect 46566 19660 46572 19672
rect 46624 19660 46630 19712
rect 48958 19660 48964 19712
rect 49016 19700 49022 19712
rect 49513 19703 49571 19709
rect 49513 19700 49525 19703
rect 49016 19672 49525 19700
rect 49016 19660 49022 19672
rect 49513 19669 49525 19672
rect 49559 19669 49571 19703
rect 49513 19663 49571 19669
rect 51721 19703 51779 19709
rect 51721 19669 51733 19703
rect 51767 19700 51779 19703
rect 51810 19700 51816 19712
rect 51767 19672 51816 19700
rect 51767 19669 51779 19672
rect 51721 19663 51779 19669
rect 51810 19660 51816 19672
rect 51868 19660 51874 19712
rect 51920 19700 51948 19799
rect 52086 19796 52092 19808
rect 52144 19796 52150 19848
rect 52181 19839 52239 19845
rect 52181 19805 52193 19839
rect 52227 19805 52239 19839
rect 52181 19799 52239 19805
rect 52917 19839 52975 19845
rect 52917 19805 52929 19839
rect 52963 19836 52975 19839
rect 53098 19836 53104 19848
rect 52963 19808 53104 19836
rect 52963 19805 52975 19808
rect 52917 19799 52975 19805
rect 52196 19768 52224 19799
rect 53098 19796 53104 19808
rect 53156 19836 53162 19848
rect 53650 19836 53656 19848
rect 53156 19808 53656 19836
rect 53156 19796 53162 19808
rect 53650 19796 53656 19808
rect 53708 19796 53714 19848
rect 53742 19796 53748 19848
rect 53800 19836 53806 19848
rect 53800 19808 53845 19836
rect 53800 19796 53806 19808
rect 54754 19796 54760 19848
rect 54812 19836 54818 19848
rect 55508 19845 55536 19944
rect 55582 19864 55588 19916
rect 55640 19904 55646 19916
rect 56318 19904 56324 19916
rect 55640 19876 56324 19904
rect 55640 19864 55646 19876
rect 56318 19864 56324 19876
rect 56376 19864 56382 19916
rect 55493 19839 55551 19845
rect 55493 19836 55505 19839
rect 54812 19808 55505 19836
rect 54812 19796 54818 19808
rect 55493 19805 55505 19808
rect 55539 19805 55551 19839
rect 55493 19799 55551 19805
rect 53834 19768 53840 19780
rect 52196 19740 53840 19768
rect 53834 19728 53840 19740
rect 53892 19728 53898 19780
rect 56597 19771 56655 19777
rect 56597 19737 56609 19771
rect 56643 19737 56655 19771
rect 56597 19731 56655 19737
rect 52454 19700 52460 19712
rect 51920 19672 52460 19700
rect 52454 19660 52460 19672
rect 52512 19660 52518 19712
rect 53282 19700 53288 19712
rect 53243 19672 53288 19700
rect 53282 19660 53288 19672
rect 53340 19660 53346 19712
rect 55861 19703 55919 19709
rect 55861 19669 55873 19703
rect 55907 19700 55919 19703
rect 56612 19700 56640 19731
rect 57330 19728 57336 19780
rect 57388 19728 57394 19780
rect 55907 19672 56640 19700
rect 55907 19669 55919 19672
rect 55861 19663 55919 19669
rect 1104 19610 58880 19632
rect 1104 19558 15398 19610
rect 15450 19558 15462 19610
rect 15514 19558 15526 19610
rect 15578 19558 15590 19610
rect 15642 19558 15654 19610
rect 15706 19558 29846 19610
rect 29898 19558 29910 19610
rect 29962 19558 29974 19610
rect 30026 19558 30038 19610
rect 30090 19558 30102 19610
rect 30154 19558 44294 19610
rect 44346 19558 44358 19610
rect 44410 19558 44422 19610
rect 44474 19558 44486 19610
rect 44538 19558 44550 19610
rect 44602 19558 58880 19610
rect 1104 19536 58880 19558
rect 5261 19499 5319 19505
rect 5261 19465 5273 19499
rect 5307 19496 5319 19499
rect 6178 19496 6184 19508
rect 5307 19468 6184 19496
rect 5307 19465 5319 19468
rect 5261 19459 5319 19465
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 7377 19499 7435 19505
rect 7377 19465 7389 19499
rect 7423 19496 7435 19499
rect 7423 19468 7880 19496
rect 7423 19465 7435 19468
rect 7377 19459 7435 19465
rect 4246 19388 4252 19440
rect 4304 19388 4310 19440
rect 5350 19388 5356 19440
rect 5408 19428 5414 19440
rect 7650 19428 7656 19440
rect 5408 19400 7656 19428
rect 5408 19388 5414 19400
rect 7650 19388 7656 19400
rect 7708 19388 7714 19440
rect 7852 19437 7880 19468
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 9732 19468 10241 19496
rect 9732 19456 9738 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 10229 19459 10287 19465
rect 10873 19499 10931 19505
rect 10873 19465 10885 19499
rect 10919 19496 10931 19499
rect 11330 19496 11336 19508
rect 10919 19468 11336 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 11330 19456 11336 19468
rect 11388 19456 11394 19508
rect 12437 19499 12495 19505
rect 12437 19465 12449 19499
rect 12483 19496 12495 19499
rect 12526 19496 12532 19508
rect 12483 19468 12532 19496
rect 12483 19465 12495 19468
rect 12437 19459 12495 19465
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 13998 19456 14004 19508
rect 14056 19496 14062 19508
rect 14277 19499 14335 19505
rect 14277 19496 14289 19499
rect 14056 19468 14289 19496
rect 14056 19456 14062 19468
rect 14277 19465 14289 19468
rect 14323 19465 14335 19499
rect 14277 19459 14335 19465
rect 14366 19456 14372 19508
rect 14424 19496 14430 19508
rect 16761 19499 16819 19505
rect 16761 19496 16773 19499
rect 14424 19468 16773 19496
rect 14424 19456 14430 19468
rect 16761 19465 16773 19468
rect 16807 19496 16819 19499
rect 17402 19496 17408 19508
rect 16807 19468 17408 19496
rect 16807 19465 16819 19468
rect 16761 19459 16819 19465
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 18693 19499 18751 19505
rect 18693 19465 18705 19499
rect 18739 19496 18751 19499
rect 18782 19496 18788 19508
rect 18739 19468 18788 19496
rect 18739 19465 18751 19468
rect 18693 19459 18751 19465
rect 18782 19456 18788 19468
rect 18840 19496 18846 19508
rect 19702 19496 19708 19508
rect 18840 19468 19708 19496
rect 18840 19456 18846 19468
rect 19702 19456 19708 19468
rect 19760 19456 19766 19508
rect 23382 19496 23388 19508
rect 22572 19468 23388 19496
rect 7837 19431 7895 19437
rect 7837 19397 7849 19431
rect 7883 19397 7895 19431
rect 11422 19428 11428 19440
rect 7837 19391 7895 19397
rect 10980 19400 11428 19428
rect 2130 19360 2136 19372
rect 2091 19332 2136 19360
rect 2130 19320 2136 19332
rect 2188 19320 2194 19372
rect 6362 19320 6368 19372
rect 6420 19360 6426 19372
rect 6549 19363 6607 19369
rect 6549 19360 6561 19363
rect 6420 19332 6561 19360
rect 6420 19320 6426 19332
rect 6549 19329 6561 19332
rect 6595 19329 6607 19363
rect 6549 19323 6607 19329
rect 6641 19363 6699 19369
rect 6641 19329 6653 19363
rect 6687 19360 6699 19363
rect 7098 19360 7104 19372
rect 6687 19332 7104 19360
rect 6687 19329 6699 19332
rect 6641 19323 6699 19329
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 7193 19363 7251 19369
rect 7193 19329 7205 19363
rect 7239 19360 7251 19363
rect 10226 19360 10232 19372
rect 7239 19332 10232 19360
rect 7239 19329 7251 19332
rect 7193 19323 7251 19329
rect 10226 19320 10232 19332
rect 10284 19320 10290 19372
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10870 19360 10876 19372
rect 10367 19332 10876 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 10980 19369 11008 19400
rect 11422 19388 11428 19400
rect 11480 19428 11486 19440
rect 12342 19428 12348 19440
rect 11480 19400 12348 19428
rect 11480 19388 11486 19400
rect 12342 19388 12348 19400
rect 12400 19388 12406 19440
rect 14016 19428 14044 19456
rect 18230 19428 18236 19440
rect 12544 19400 14044 19428
rect 17420 19400 18236 19428
rect 10965 19363 11023 19369
rect 10965 19329 10977 19363
rect 11011 19329 11023 19363
rect 11698 19360 11704 19372
rect 11659 19332 11704 19360
rect 10965 19323 11023 19329
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19360 11851 19363
rect 11882 19360 11888 19372
rect 11839 19332 11888 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 12544 19369 12572 19400
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19329 12587 19363
rect 12986 19360 12992 19372
rect 12947 19332 12992 19360
rect 12529 19323 12587 19329
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 17420 19369 17448 19400
rect 18230 19388 18236 19400
rect 18288 19388 18294 19440
rect 19334 19388 19340 19440
rect 19392 19428 19398 19440
rect 21913 19431 21971 19437
rect 21913 19428 21925 19431
rect 19392 19400 21925 19428
rect 19392 19388 19398 19400
rect 21913 19397 21925 19400
rect 21959 19397 21971 19431
rect 22572 19428 22600 19468
rect 23382 19456 23388 19468
rect 23440 19456 23446 19508
rect 23474 19456 23480 19508
rect 23532 19496 23538 19508
rect 24765 19499 24823 19505
rect 24765 19496 24777 19499
rect 23532 19468 24777 19496
rect 23532 19456 23538 19468
rect 24765 19465 24777 19468
rect 24811 19465 24823 19499
rect 26421 19499 26479 19505
rect 26421 19496 26433 19499
rect 24765 19459 24823 19465
rect 26206 19468 26433 19496
rect 25130 19428 25136 19440
rect 21913 19391 21971 19397
rect 22480 19400 22600 19428
rect 23966 19400 25136 19428
rect 17405 19363 17463 19369
rect 15068 19332 17356 19360
rect 15068 19320 15074 19332
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 3513 19295 3571 19301
rect 3513 19292 3525 19295
rect 2516 19264 3525 19292
rect 2516 19233 2544 19264
rect 3513 19261 3525 19264
rect 3559 19261 3571 19295
rect 3513 19255 3571 19261
rect 3789 19295 3847 19301
rect 3789 19261 3801 19295
rect 3835 19292 3847 19295
rect 3878 19292 3884 19304
rect 3835 19264 3884 19292
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 4246 19252 4252 19304
rect 4304 19292 4310 19304
rect 6914 19292 6920 19304
rect 4304 19264 6920 19292
rect 4304 19252 4310 19264
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 7024 19264 12434 19292
rect 2501 19227 2559 19233
rect 2501 19193 2513 19227
rect 2547 19193 2559 19227
rect 2501 19187 2559 19193
rect 5442 19184 5448 19236
rect 5500 19224 5506 19236
rect 7024 19224 7052 19264
rect 9122 19224 9128 19236
rect 5500 19196 7052 19224
rect 9083 19196 9128 19224
rect 5500 19184 5506 19196
rect 9122 19184 9128 19196
rect 9180 19184 9186 19236
rect 12406 19224 12434 19264
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 13262 19292 13268 19304
rect 12952 19264 13268 19292
rect 12952 19252 12958 19264
rect 13262 19252 13268 19264
rect 13320 19252 13326 19304
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16025 19295 16083 19301
rect 16025 19292 16037 19295
rect 15611 19264 16037 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 16025 19261 16037 19264
rect 16071 19292 16083 19295
rect 17034 19292 17040 19304
rect 16071 19264 17040 19292
rect 16071 19261 16083 19264
rect 16025 19255 16083 19261
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 17328 19292 17356 19332
rect 17405 19329 17417 19363
rect 17451 19329 17463 19363
rect 17865 19363 17923 19369
rect 17865 19360 17877 19363
rect 17405 19323 17463 19329
rect 17512 19332 17877 19360
rect 17512 19292 17540 19332
rect 17865 19329 17877 19332
rect 17911 19329 17923 19363
rect 17865 19323 17923 19329
rect 17954 19320 17960 19372
rect 18012 19360 18018 19372
rect 18509 19363 18567 19369
rect 18012 19332 18057 19360
rect 18012 19320 18018 19332
rect 18509 19329 18521 19363
rect 18555 19360 18567 19363
rect 18874 19360 18880 19372
rect 18555 19332 18880 19360
rect 18555 19329 18567 19332
rect 18509 19323 18567 19329
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19978 19360 19984 19372
rect 19939 19332 19984 19360
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19360 22063 19363
rect 22370 19360 22376 19372
rect 22051 19332 22376 19360
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 22480 19369 22508 19400
rect 25130 19388 25136 19400
rect 25188 19388 25194 19440
rect 22465 19363 22523 19369
rect 22465 19329 22477 19363
rect 22511 19329 22523 19363
rect 24854 19360 24860 19372
rect 24815 19332 24860 19360
rect 22465 19323 22523 19329
rect 24854 19320 24860 19332
rect 24912 19320 24918 19372
rect 25501 19363 25559 19369
rect 25501 19329 25513 19363
rect 25547 19360 25559 19363
rect 26206 19360 26234 19468
rect 26421 19465 26433 19468
rect 26467 19496 26479 19499
rect 27798 19496 27804 19508
rect 26467 19468 27804 19496
rect 26467 19465 26479 19468
rect 26421 19459 26479 19465
rect 27798 19456 27804 19468
rect 27856 19456 27862 19508
rect 31018 19496 31024 19508
rect 30979 19468 31024 19496
rect 31018 19456 31024 19468
rect 31076 19456 31082 19508
rect 36262 19496 36268 19508
rect 31128 19468 36268 19496
rect 27246 19428 27252 19440
rect 27207 19400 27252 19428
rect 27246 19388 27252 19400
rect 27304 19388 27310 19440
rect 28905 19431 28963 19437
rect 28905 19397 28917 19431
rect 28951 19428 28963 19431
rect 30558 19428 30564 19440
rect 28951 19400 30564 19428
rect 28951 19397 28963 19400
rect 28905 19391 28963 19397
rect 30558 19388 30564 19400
rect 30616 19388 30622 19440
rect 25547 19332 26234 19360
rect 25547 19329 25559 19332
rect 25501 19323 25559 19329
rect 17328 19264 17540 19292
rect 19610 19252 19616 19304
rect 19668 19292 19674 19304
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 19668 19264 19901 19292
rect 19668 19252 19674 19264
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 22741 19295 22799 19301
rect 22741 19292 22753 19295
rect 19889 19255 19947 19261
rect 22066 19264 22753 19292
rect 16758 19224 16764 19236
rect 12406 19196 16764 19224
rect 16758 19184 16764 19196
rect 16816 19224 16822 19236
rect 19337 19227 19395 19233
rect 19337 19224 19349 19227
rect 16816 19196 19349 19224
rect 16816 19184 16822 19196
rect 19337 19193 19349 19196
rect 19383 19224 19395 19227
rect 19426 19224 19432 19236
rect 19383 19196 19432 19224
rect 19383 19193 19395 19196
rect 19337 19187 19395 19193
rect 19426 19184 19432 19196
rect 19484 19184 19490 19236
rect 20349 19227 20407 19233
rect 20349 19193 20361 19227
rect 20395 19224 20407 19227
rect 22066 19224 22094 19264
rect 22741 19261 22753 19264
rect 22787 19261 22799 19295
rect 22741 19255 22799 19261
rect 25038 19252 25044 19304
rect 25096 19292 25102 19304
rect 25409 19295 25467 19301
rect 25409 19292 25421 19295
rect 25096 19264 25421 19292
rect 25096 19252 25102 19264
rect 25409 19261 25421 19264
rect 25455 19261 25467 19295
rect 25409 19255 25467 19261
rect 20395 19196 22094 19224
rect 20395 19193 20407 19196
rect 20349 19187 20407 19193
rect 23750 19184 23756 19236
rect 23808 19224 23814 19236
rect 26206 19224 26234 19332
rect 27065 19363 27123 19369
rect 27065 19329 27077 19363
rect 27111 19329 27123 19363
rect 31018 19360 31024 19372
rect 27065 19323 27123 19329
rect 28460 19332 31024 19360
rect 27080 19292 27108 19323
rect 28460 19292 28488 19332
rect 31018 19320 31024 19332
rect 31076 19320 31082 19372
rect 31128 19369 31156 19468
rect 36262 19456 36268 19468
rect 36320 19456 36326 19508
rect 40310 19456 40316 19508
rect 40368 19496 40374 19508
rect 40957 19499 41015 19505
rect 40957 19496 40969 19499
rect 40368 19468 40969 19496
rect 40368 19456 40374 19468
rect 40957 19465 40969 19468
rect 41003 19465 41015 19499
rect 40957 19459 41015 19465
rect 42150 19456 42156 19508
rect 42208 19496 42214 19508
rect 42521 19499 42579 19505
rect 42521 19496 42533 19499
rect 42208 19468 42533 19496
rect 42208 19456 42214 19468
rect 42521 19465 42533 19468
rect 42567 19465 42579 19499
rect 43254 19496 43260 19508
rect 43215 19468 43260 19496
rect 42521 19459 42579 19465
rect 43254 19456 43260 19468
rect 43312 19456 43318 19508
rect 48314 19456 48320 19508
rect 48372 19496 48378 19508
rect 48593 19499 48651 19505
rect 48593 19496 48605 19499
rect 48372 19468 48605 19496
rect 48372 19456 48378 19468
rect 48593 19465 48605 19468
rect 48639 19465 48651 19499
rect 48593 19459 48651 19465
rect 51350 19456 51356 19508
rect 51408 19496 51414 19508
rect 51629 19499 51687 19505
rect 51629 19496 51641 19499
rect 51408 19468 51641 19496
rect 51408 19456 51414 19468
rect 51629 19465 51641 19468
rect 51675 19465 51687 19499
rect 51629 19459 51687 19465
rect 53006 19456 53012 19508
rect 53064 19496 53070 19508
rect 53193 19499 53251 19505
rect 53193 19496 53205 19499
rect 53064 19468 53205 19496
rect 53064 19456 53070 19468
rect 53193 19465 53205 19468
rect 53239 19465 53251 19499
rect 53650 19496 53656 19508
rect 53563 19468 53656 19496
rect 53193 19459 53251 19465
rect 53650 19456 53656 19468
rect 53708 19496 53714 19508
rect 56045 19499 56103 19505
rect 56045 19496 56057 19499
rect 53708 19468 56057 19496
rect 53708 19456 53714 19468
rect 56045 19465 56057 19468
rect 56091 19465 56103 19499
rect 56045 19459 56103 19465
rect 35342 19428 35348 19440
rect 33626 19400 35348 19428
rect 35342 19388 35348 19400
rect 35400 19388 35406 19440
rect 41046 19428 41052 19440
rect 40710 19400 41052 19428
rect 41046 19388 41052 19400
rect 41104 19388 41110 19440
rect 31113 19363 31171 19369
rect 31113 19329 31125 19363
rect 31159 19329 31171 19363
rect 32125 19363 32183 19369
rect 32125 19360 32137 19363
rect 31113 19323 31171 19329
rect 31220 19332 32137 19360
rect 29454 19292 29460 19304
rect 27080 19264 28488 19292
rect 29367 19264 29460 19292
rect 29454 19252 29460 19264
rect 29512 19292 29518 19304
rect 30190 19292 30196 19304
rect 29512 19264 30196 19292
rect 29512 19252 29518 19264
rect 30190 19252 30196 19264
rect 30248 19252 30254 19304
rect 31220 19292 31248 19332
rect 32125 19329 32137 19332
rect 32171 19329 32183 19363
rect 34606 19360 34612 19372
rect 34567 19332 34612 19360
rect 32125 19323 32183 19329
rect 34606 19320 34612 19332
rect 34664 19320 34670 19372
rect 35250 19320 35256 19372
rect 35308 19360 35314 19372
rect 36173 19363 36231 19369
rect 36173 19360 36185 19363
rect 35308 19332 36185 19360
rect 35308 19320 35314 19332
rect 36173 19329 36185 19332
rect 36219 19329 36231 19363
rect 36173 19323 36231 19329
rect 37458 19320 37464 19372
rect 37516 19360 37522 19372
rect 37553 19363 37611 19369
rect 37553 19360 37565 19363
rect 37516 19332 37565 19360
rect 37516 19320 37522 19332
rect 37553 19329 37565 19332
rect 37599 19329 37611 19363
rect 39206 19360 39212 19372
rect 39167 19332 39212 19360
rect 37553 19323 37611 19329
rect 39206 19320 39212 19332
rect 39264 19320 39270 19372
rect 41598 19360 41604 19372
rect 41559 19332 41604 19360
rect 41598 19320 41604 19332
rect 41656 19320 41662 19372
rect 42610 19360 42616 19372
rect 42571 19332 42616 19360
rect 42610 19320 42616 19332
rect 42668 19320 42674 19372
rect 43070 19360 43076 19372
rect 43031 19332 43076 19360
rect 43070 19320 43076 19332
rect 43128 19320 43134 19372
rect 43272 19360 43300 19456
rect 46566 19428 46572 19440
rect 44468 19400 45692 19428
rect 46527 19400 46572 19428
rect 43717 19363 43775 19369
rect 43717 19360 43729 19363
rect 43272 19332 43729 19360
rect 43717 19329 43729 19332
rect 43763 19329 43775 19363
rect 43990 19360 43996 19372
rect 43903 19332 43996 19360
rect 43717 19323 43775 19329
rect 43990 19320 43996 19332
rect 44048 19360 44054 19372
rect 44468 19360 44496 19400
rect 44634 19360 44640 19372
rect 44048 19332 44496 19360
rect 44595 19332 44640 19360
rect 44048 19320 44054 19332
rect 44634 19320 44640 19332
rect 44692 19320 44698 19372
rect 45370 19360 45376 19372
rect 45331 19332 45376 19360
rect 45370 19320 45376 19332
rect 45428 19320 45434 19372
rect 45664 19369 45692 19400
rect 46566 19388 46572 19400
rect 46624 19388 46630 19440
rect 50338 19428 50344 19440
rect 49344 19400 50344 19428
rect 45649 19363 45707 19369
rect 45649 19329 45661 19363
rect 45695 19360 45707 19363
rect 45738 19360 45744 19372
rect 45695 19332 45744 19360
rect 45695 19329 45707 19332
rect 45649 19323 45707 19329
rect 45738 19320 45744 19332
rect 45796 19360 45802 19372
rect 46290 19360 46296 19372
rect 45796 19332 46060 19360
rect 46251 19332 46296 19360
rect 45796 19320 45802 19332
rect 30392 19264 31248 19292
rect 32401 19295 32459 19301
rect 26602 19224 26608 19236
rect 23808 19196 26608 19224
rect 23808 19184 23814 19196
rect 26602 19184 26608 19196
rect 26660 19184 26666 19236
rect 30392 19168 30420 19264
rect 32401 19261 32413 19295
rect 32447 19292 32459 19295
rect 32490 19292 32496 19304
rect 32447 19264 32496 19292
rect 32447 19261 32459 19264
rect 32401 19255 32459 19261
rect 32490 19252 32496 19264
rect 32548 19252 32554 19304
rect 34517 19295 34575 19301
rect 34517 19292 34529 19295
rect 33888 19264 34529 19292
rect 33888 19168 33916 19264
rect 34517 19261 34529 19264
rect 34563 19261 34575 19295
rect 35434 19292 35440 19304
rect 35395 19264 35440 19292
rect 34517 19255 34575 19261
rect 35434 19252 35440 19264
rect 35492 19252 35498 19304
rect 35897 19295 35955 19301
rect 35897 19261 35909 19295
rect 35943 19292 35955 19295
rect 36078 19292 36084 19304
rect 35943 19264 36084 19292
rect 35943 19261 35955 19264
rect 35897 19255 35955 19261
rect 36078 19252 36084 19264
rect 36136 19252 36142 19304
rect 37645 19295 37703 19301
rect 37645 19261 37657 19295
rect 37691 19261 37703 19295
rect 38378 19292 38384 19304
rect 38339 19264 38384 19292
rect 37645 19255 37703 19261
rect 35066 19184 35072 19236
rect 35124 19224 35130 19236
rect 37660 19224 37688 19255
rect 38378 19252 38384 19264
rect 38436 19252 38442 19304
rect 39485 19295 39543 19301
rect 39485 19261 39497 19295
rect 39531 19292 39543 19295
rect 41417 19295 41475 19301
rect 41417 19292 41429 19295
rect 39531 19264 41429 19292
rect 39531 19261 39543 19264
rect 39485 19255 39543 19261
rect 41417 19261 41429 19264
rect 41463 19261 41475 19295
rect 46032 19292 46060 19332
rect 46290 19320 46296 19332
rect 46348 19320 46354 19372
rect 47946 19360 47952 19372
rect 47907 19332 47952 19360
rect 47946 19320 47952 19332
rect 48004 19320 48010 19372
rect 48866 19360 48872 19372
rect 48827 19332 48872 19360
rect 48866 19320 48872 19332
rect 48924 19320 48930 19372
rect 49344 19369 49372 19400
rect 50338 19388 50344 19400
rect 50396 19388 50402 19440
rect 50798 19388 50804 19440
rect 50856 19428 50862 19440
rect 50856 19400 53604 19428
rect 50856 19388 50862 19400
rect 49329 19363 49387 19369
rect 49329 19329 49341 19363
rect 49375 19329 49387 19363
rect 49329 19323 49387 19329
rect 51074 19320 51080 19372
rect 51132 19360 51138 19372
rect 51629 19363 51687 19369
rect 51629 19360 51641 19363
rect 51132 19332 51641 19360
rect 51132 19320 51138 19332
rect 51629 19329 51641 19332
rect 51675 19329 51687 19363
rect 51810 19360 51816 19372
rect 51771 19332 51816 19360
rect 51629 19323 51687 19329
rect 51810 19320 51816 19332
rect 51868 19320 51874 19372
rect 52748 19369 52776 19400
rect 52733 19363 52791 19369
rect 52733 19329 52745 19363
rect 52779 19329 52791 19363
rect 52733 19323 52791 19329
rect 52822 19320 52828 19372
rect 52880 19360 52886 19372
rect 52880 19332 52925 19360
rect 52880 19320 52886 19332
rect 53006 19320 53012 19372
rect 53064 19360 53070 19372
rect 53064 19332 53109 19360
rect 53064 19320 53070 19332
rect 46474 19292 46480 19304
rect 46032 19264 46480 19292
rect 41417 19255 41475 19261
rect 46474 19252 46480 19264
rect 46532 19252 46538 19304
rect 47581 19295 47639 19301
rect 47581 19261 47593 19295
rect 47627 19292 47639 19295
rect 47670 19292 47676 19304
rect 47627 19264 47676 19292
rect 47627 19261 47639 19264
rect 47581 19255 47639 19261
rect 47670 19252 47676 19264
rect 47728 19252 47734 19304
rect 48038 19292 48044 19304
rect 47999 19264 48044 19292
rect 48038 19252 48044 19264
rect 48096 19252 48102 19304
rect 48593 19295 48651 19301
rect 48593 19261 48605 19295
rect 48639 19261 48651 19295
rect 48593 19255 48651 19261
rect 48777 19295 48835 19301
rect 48777 19261 48789 19295
rect 48823 19292 48835 19295
rect 48958 19292 48964 19304
rect 48823 19264 48964 19292
rect 48823 19261 48835 19264
rect 48777 19255 48835 19261
rect 35124 19196 37688 19224
rect 48608 19224 48636 19255
rect 48958 19252 48964 19264
rect 49016 19252 49022 19304
rect 49510 19292 49516 19304
rect 49471 19264 49516 19292
rect 49510 19252 49516 19264
rect 49568 19252 49574 19304
rect 51166 19292 51172 19304
rect 51127 19264 51172 19292
rect 51166 19252 51172 19264
rect 51224 19252 51230 19304
rect 53576 19292 53604 19400
rect 53668 19369 53696 19456
rect 57330 19428 57336 19440
rect 55798 19400 57336 19428
rect 57330 19388 57336 19400
rect 57388 19388 57394 19440
rect 53653 19363 53711 19369
rect 53653 19329 53665 19363
rect 53699 19329 53711 19363
rect 53837 19363 53895 19369
rect 53837 19360 53849 19363
rect 53653 19323 53711 19329
rect 53760 19332 53849 19360
rect 53760 19292 53788 19332
rect 53837 19329 53849 19332
rect 53883 19360 53895 19363
rect 53926 19360 53932 19372
rect 53883 19332 53932 19360
rect 53883 19329 53895 19332
rect 53837 19323 53895 19329
rect 53926 19320 53932 19332
rect 53984 19320 53990 19372
rect 54294 19360 54300 19372
rect 54255 19332 54300 19360
rect 54294 19320 54300 19332
rect 54352 19320 54358 19372
rect 54573 19295 54631 19301
rect 54573 19292 54585 19295
rect 53576 19264 53788 19292
rect 54404 19264 54585 19292
rect 52546 19224 52552 19236
rect 48608 19196 52552 19224
rect 35124 19184 35130 19196
rect 52546 19184 52552 19196
rect 52604 19184 52610 19236
rect 53282 19184 53288 19236
rect 53340 19224 53346 19236
rect 54404 19224 54432 19264
rect 54573 19261 54585 19264
rect 54619 19261 54631 19295
rect 54573 19255 54631 19261
rect 53340 19196 54432 19224
rect 53340 19184 53346 19196
rect 3053 19159 3111 19165
rect 3053 19125 3065 19159
rect 3099 19156 3111 19159
rect 3970 19156 3976 19168
rect 3099 19128 3976 19156
rect 3099 19125 3111 19128
rect 3053 19119 3111 19125
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 5813 19159 5871 19165
rect 5813 19125 5825 19159
rect 5859 19156 5871 19159
rect 9582 19156 9588 19168
rect 5859 19128 9588 19156
rect 5859 19125 5871 19128
rect 5813 19119 5871 19125
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 11330 19116 11336 19168
rect 11388 19156 11394 19168
rect 13170 19156 13176 19168
rect 11388 19128 13176 19156
rect 11388 19116 11394 19128
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 17310 19156 17316 19168
rect 17271 19128 17316 19156
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 21174 19156 21180 19168
rect 21135 19128 21180 19156
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 24210 19156 24216 19168
rect 24171 19128 24216 19156
rect 24210 19116 24216 19128
rect 24268 19116 24274 19168
rect 25777 19159 25835 19165
rect 25777 19125 25789 19159
rect 25823 19156 25835 19159
rect 26142 19156 26148 19168
rect 25823 19128 26148 19156
rect 25823 19125 25835 19128
rect 25777 19119 25835 19125
rect 26142 19116 26148 19128
rect 26200 19116 26206 19168
rect 30374 19156 30380 19168
rect 30335 19128 30380 19156
rect 30374 19116 30380 19128
rect 30432 19116 30438 19168
rect 33870 19156 33876 19168
rect 33831 19128 33876 19156
rect 33870 19116 33876 19128
rect 33928 19116 33934 19168
rect 44634 19116 44640 19168
rect 44692 19156 44698 19168
rect 44821 19159 44879 19165
rect 44821 19156 44833 19159
rect 44692 19128 44833 19156
rect 44692 19116 44698 19128
rect 44821 19125 44833 19128
rect 44867 19125 44879 19159
rect 44821 19119 44879 19125
rect 46474 19116 46480 19168
rect 46532 19156 46538 19168
rect 51166 19156 51172 19168
rect 46532 19128 51172 19156
rect 46532 19116 46538 19128
rect 51166 19116 51172 19128
rect 51224 19116 51230 19168
rect 53834 19156 53840 19168
rect 53795 19128 53840 19156
rect 53834 19116 53840 19128
rect 53892 19116 53898 19168
rect 1104 19066 58880 19088
rect 1104 19014 8174 19066
rect 8226 19014 8238 19066
rect 8290 19014 8302 19066
rect 8354 19014 8366 19066
rect 8418 19014 8430 19066
rect 8482 19014 22622 19066
rect 22674 19014 22686 19066
rect 22738 19014 22750 19066
rect 22802 19014 22814 19066
rect 22866 19014 22878 19066
rect 22930 19014 37070 19066
rect 37122 19014 37134 19066
rect 37186 19014 37198 19066
rect 37250 19014 37262 19066
rect 37314 19014 37326 19066
rect 37378 19014 51518 19066
rect 51570 19014 51582 19066
rect 51634 19014 51646 19066
rect 51698 19014 51710 19066
rect 51762 19014 51774 19066
rect 51826 19014 58880 19066
rect 1104 18992 58880 19014
rect 9585 18955 9643 18961
rect 9585 18921 9597 18955
rect 9631 18952 9643 18955
rect 11790 18952 11796 18964
rect 9631 18924 11796 18952
rect 9631 18921 9643 18924
rect 9585 18915 9643 18921
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 11900 18924 14412 18952
rect 3145 18887 3203 18893
rect 3145 18853 3157 18887
rect 3191 18853 3203 18887
rect 11330 18884 11336 18896
rect 3145 18847 3203 18853
rect 10336 18856 11336 18884
rect 2222 18816 2228 18828
rect 2135 18788 2228 18816
rect 2222 18776 2228 18788
rect 2280 18816 2286 18828
rect 3160 18816 3188 18847
rect 3973 18819 4031 18825
rect 3973 18816 3985 18819
rect 2280 18788 3985 18816
rect 2280 18776 2286 18788
rect 3973 18785 3985 18788
rect 4019 18785 4031 18819
rect 3973 18779 4031 18785
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18748 3019 18751
rect 3050 18748 3056 18760
rect 3007 18720 3056 18748
rect 3007 18717 3019 18720
rect 2961 18711 3019 18717
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 4246 18748 4252 18760
rect 4207 18720 4252 18748
rect 4246 18708 4252 18720
rect 4304 18708 4310 18760
rect 5902 18748 5908 18760
rect 5863 18720 5908 18748
rect 5902 18708 5908 18720
rect 5960 18708 5966 18760
rect 10336 18757 10364 18856
rect 11330 18844 11336 18856
rect 11388 18844 11394 18896
rect 11514 18844 11520 18896
rect 11572 18884 11578 18896
rect 11900 18884 11928 18924
rect 11572 18856 11928 18884
rect 11572 18844 11578 18856
rect 10873 18819 10931 18825
rect 10873 18785 10885 18819
rect 10919 18816 10931 18819
rect 12989 18819 13047 18825
rect 12989 18816 13001 18819
rect 10919 18788 13001 18816
rect 10919 18785 10931 18788
rect 10873 18779 10931 18785
rect 12989 18785 13001 18788
rect 13035 18785 13047 18819
rect 12989 18779 13047 18785
rect 13354 18776 13360 18828
rect 13412 18816 13418 18828
rect 14277 18819 14335 18825
rect 14277 18816 14289 18819
rect 13412 18788 14289 18816
rect 13412 18776 13418 18788
rect 14277 18785 14289 18788
rect 14323 18785 14335 18819
rect 14277 18779 14335 18785
rect 6365 18751 6423 18757
rect 6365 18717 6377 18751
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 9677 18751 9735 18757
rect 9677 18717 9689 18751
rect 9723 18748 9735 18751
rect 10321 18751 10379 18757
rect 9723 18720 10272 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 6380 18680 6408 18711
rect 6638 18680 6644 18692
rect 2516 18652 6408 18680
rect 6599 18652 6644 18680
rect 2516 18621 2544 18652
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 7098 18640 7104 18692
rect 7156 18640 7162 18692
rect 9033 18683 9091 18689
rect 9033 18649 9045 18683
rect 9079 18680 9091 18683
rect 9858 18680 9864 18692
rect 9079 18652 9864 18680
rect 9079 18649 9091 18652
rect 9033 18643 9091 18649
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 10244 18680 10272 18720
rect 10321 18717 10333 18751
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18748 11023 18751
rect 11011 18720 11744 18748
rect 11011 18717 11023 18720
rect 10965 18711 11023 18717
rect 10244 18652 10916 18680
rect 2501 18615 2559 18621
rect 2501 18581 2513 18615
rect 2547 18581 2559 18615
rect 4890 18612 4896 18624
rect 4851 18584 4896 18612
rect 2501 18575 2559 18581
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 5813 18615 5871 18621
rect 5813 18581 5825 18615
rect 5859 18612 5871 18615
rect 7282 18612 7288 18624
rect 5859 18584 7288 18612
rect 5859 18581 5871 18584
rect 5813 18575 5871 18581
rect 7282 18572 7288 18584
rect 7340 18572 7346 18624
rect 7466 18572 7472 18624
rect 7524 18612 7530 18624
rect 8113 18615 8171 18621
rect 8113 18612 8125 18615
rect 7524 18584 8125 18612
rect 7524 18572 7530 18584
rect 8113 18581 8125 18584
rect 8159 18581 8171 18615
rect 10226 18612 10232 18624
rect 10187 18584 10232 18612
rect 8113 18575 8171 18581
rect 10226 18572 10232 18584
rect 10284 18572 10290 18624
rect 10888 18612 10916 18652
rect 11330 18612 11336 18624
rect 10888 18584 11336 18612
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 11514 18612 11520 18624
rect 11475 18584 11520 18612
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 11716 18612 11744 18720
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 14384 18757 14412 18924
rect 14844 18924 18736 18952
rect 14369 18751 14427 18757
rect 13320 18720 13365 18748
rect 13320 18708 13326 18720
rect 14369 18717 14381 18751
rect 14415 18717 14427 18751
rect 14369 18711 14427 18717
rect 13722 18640 13728 18692
rect 13780 18680 13786 18692
rect 14844 18680 14872 18924
rect 15102 18816 15108 18828
rect 15063 18788 15108 18816
rect 15102 18776 15108 18788
rect 15160 18776 15166 18828
rect 16301 18819 16359 18825
rect 16301 18785 16313 18819
rect 16347 18816 16359 18819
rect 18598 18816 18604 18828
rect 16347 18788 18604 18816
rect 16347 18785 16359 18788
rect 16301 18779 16359 18785
rect 18598 18776 18604 18788
rect 18656 18776 18662 18828
rect 18708 18816 18736 18924
rect 20990 18912 20996 18964
rect 21048 18952 21054 18964
rect 21085 18955 21143 18961
rect 21085 18952 21097 18955
rect 21048 18924 21097 18952
rect 21048 18912 21054 18924
rect 21085 18921 21097 18924
rect 21131 18921 21143 18955
rect 21085 18915 21143 18921
rect 22741 18955 22799 18961
rect 22741 18921 22753 18955
rect 22787 18952 22799 18955
rect 26050 18952 26056 18964
rect 22787 18924 26056 18952
rect 22787 18921 22799 18924
rect 22741 18915 22799 18921
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 28074 18912 28080 18964
rect 28132 18952 28138 18964
rect 28994 18952 29000 18964
rect 28132 18924 28580 18952
rect 28955 18924 29000 18952
rect 28132 18912 28138 18924
rect 19610 18844 19616 18896
rect 19668 18884 19674 18896
rect 20901 18887 20959 18893
rect 20901 18884 20913 18887
rect 19668 18856 20913 18884
rect 19668 18844 19674 18856
rect 20901 18853 20913 18856
rect 20947 18853 20959 18887
rect 25041 18887 25099 18893
rect 25041 18884 25053 18887
rect 20901 18847 20959 18853
rect 22066 18856 25053 18884
rect 19705 18819 19763 18825
rect 19705 18816 19717 18819
rect 18708 18788 19717 18816
rect 19705 18785 19717 18788
rect 19751 18816 19763 18819
rect 19978 18816 19984 18828
rect 19751 18788 19984 18816
rect 19751 18785 19763 18788
rect 19705 18779 19763 18785
rect 19978 18776 19984 18788
rect 20036 18816 20042 18828
rect 22066 18816 22094 18856
rect 25041 18853 25053 18856
rect 25087 18853 25099 18887
rect 28552 18884 28580 18924
rect 28994 18912 29000 18924
rect 29052 18912 29058 18964
rect 34330 18912 34336 18964
rect 34388 18952 34394 18964
rect 38746 18952 38752 18964
rect 34388 18924 36860 18952
rect 38707 18924 38752 18952
rect 34388 18912 34394 18924
rect 29549 18887 29607 18893
rect 29549 18884 29561 18887
rect 28552 18856 29561 18884
rect 25041 18847 25099 18853
rect 29549 18853 29561 18856
rect 29595 18853 29607 18887
rect 29549 18847 29607 18853
rect 22370 18816 22376 18828
rect 20036 18788 22094 18816
rect 22331 18788 22376 18816
rect 20036 18776 20042 18788
rect 22370 18776 22376 18788
rect 22428 18816 22434 18828
rect 22428 18788 23520 18816
rect 22428 18776 22434 18788
rect 16022 18748 16028 18760
rect 15983 18720 16028 18748
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 18230 18708 18236 18760
rect 18288 18748 18294 18760
rect 18325 18751 18383 18757
rect 18325 18748 18337 18751
rect 18288 18720 18337 18748
rect 18288 18708 18294 18720
rect 18325 18717 18337 18720
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 20349 18751 20407 18757
rect 18472 18720 18517 18748
rect 18472 18708 18478 18720
rect 20349 18717 20361 18751
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 13780 18652 14872 18680
rect 13780 18640 13786 18652
rect 17310 18640 17316 18692
rect 17368 18640 17374 18692
rect 17604 18652 18000 18680
rect 13354 18612 13360 18624
rect 11716 18584 13360 18612
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 14550 18572 14556 18624
rect 14608 18612 14614 18624
rect 17604 18612 17632 18652
rect 17770 18612 17776 18624
rect 14608 18584 17632 18612
rect 17731 18584 17776 18612
rect 14608 18572 14614 18584
rect 17770 18572 17776 18584
rect 17828 18572 17834 18624
rect 17972 18612 18000 18652
rect 18046 18640 18052 18692
rect 18104 18680 18110 18692
rect 20257 18683 20315 18689
rect 20257 18680 20269 18683
rect 18104 18652 20269 18680
rect 18104 18640 18110 18652
rect 20257 18649 20269 18652
rect 20303 18649 20315 18683
rect 20364 18680 20392 18711
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20772 18720 21097 18748
rect 20772 18708 20778 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 21174 18708 21180 18760
rect 21232 18748 21238 18760
rect 22462 18748 22468 18760
rect 21232 18720 21277 18748
rect 22423 18720 22468 18748
rect 21232 18708 21238 18720
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 23492 18748 23520 18788
rect 23566 18776 23572 18828
rect 23624 18816 23630 18828
rect 23845 18819 23903 18825
rect 23845 18816 23857 18819
rect 23624 18788 23857 18816
rect 23624 18776 23630 18788
rect 23845 18785 23857 18788
rect 23891 18816 23903 18819
rect 27249 18819 27307 18825
rect 27249 18816 27261 18819
rect 23891 18788 27261 18816
rect 23891 18785 23903 18788
rect 23845 18779 23903 18785
rect 27249 18785 27261 18788
rect 27295 18816 27307 18819
rect 29454 18816 29460 18828
rect 27295 18788 29460 18816
rect 27295 18785 27307 18788
rect 27249 18779 27307 18785
rect 29454 18776 29460 18788
rect 29512 18776 29518 18828
rect 36725 18819 36783 18825
rect 36725 18816 36737 18819
rect 31726 18788 36737 18816
rect 23750 18748 23756 18760
rect 23492 18720 23756 18748
rect 23750 18708 23756 18720
rect 23808 18708 23814 18760
rect 24210 18708 24216 18760
rect 24268 18748 24274 18760
rect 24857 18751 24915 18757
rect 24857 18748 24869 18751
rect 24268 18720 24869 18748
rect 24268 18708 24274 18720
rect 24857 18717 24869 18720
rect 24903 18717 24915 18751
rect 25774 18748 25780 18760
rect 25735 18720 25780 18748
rect 24857 18711 24915 18717
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 25958 18748 25964 18760
rect 25919 18720 25964 18748
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 30466 18748 30472 18760
rect 30427 18720 30472 18748
rect 30466 18708 30472 18720
rect 30524 18708 30530 18760
rect 31386 18748 31392 18760
rect 31299 18720 31392 18748
rect 31386 18708 31392 18720
rect 31444 18748 31450 18760
rect 31726 18748 31754 18788
rect 36725 18785 36737 18788
rect 36771 18785 36783 18819
rect 36832 18816 36860 18924
rect 38746 18912 38752 18924
rect 38804 18912 38810 18964
rect 48593 18955 48651 18961
rect 38856 18924 47532 18952
rect 36906 18844 36912 18896
rect 36964 18884 36970 18896
rect 38856 18884 38884 18924
rect 36964 18856 38884 18884
rect 45373 18887 45431 18893
rect 36964 18844 36970 18856
rect 45373 18853 45385 18887
rect 45419 18884 45431 18887
rect 45646 18884 45652 18896
rect 45419 18856 45652 18884
rect 45419 18853 45431 18856
rect 45373 18847 45431 18853
rect 45646 18844 45652 18856
rect 45704 18844 45710 18896
rect 37369 18819 37427 18825
rect 37369 18816 37381 18819
rect 36832 18788 37381 18816
rect 36725 18779 36783 18785
rect 37369 18785 37381 18788
rect 37415 18816 37427 18819
rect 40126 18816 40132 18828
rect 37415 18788 38792 18816
rect 40087 18788 40132 18816
rect 37415 18785 37427 18788
rect 37369 18779 37427 18785
rect 31444 18720 31754 18748
rect 33781 18751 33839 18757
rect 31444 18708 31450 18720
rect 33781 18717 33793 18751
rect 33827 18717 33839 18751
rect 33781 18711 33839 18717
rect 20364 18652 21312 18680
rect 20257 18643 20315 18649
rect 21174 18612 21180 18624
rect 17972 18584 21180 18612
rect 21174 18572 21180 18584
rect 21232 18572 21238 18624
rect 21284 18612 21312 18652
rect 21358 18640 21364 18692
rect 21416 18680 21422 18692
rect 21416 18652 21461 18680
rect 21416 18640 21422 18652
rect 26142 18640 26148 18692
rect 26200 18680 26206 18692
rect 27525 18683 27583 18689
rect 27525 18680 27537 18683
rect 26200 18652 27537 18680
rect 26200 18640 26206 18652
rect 27525 18649 27537 18652
rect 27571 18649 27583 18683
rect 27525 18643 27583 18649
rect 27614 18640 27620 18692
rect 27672 18680 27678 18692
rect 27982 18680 27988 18692
rect 27672 18652 27988 18680
rect 27672 18640 27678 18652
rect 27982 18640 27988 18652
rect 28040 18640 28046 18692
rect 31941 18683 31999 18689
rect 31941 18649 31953 18683
rect 31987 18680 31999 18683
rect 32030 18680 32036 18692
rect 31987 18652 32036 18680
rect 31987 18649 31999 18652
rect 31941 18643 31999 18649
rect 32030 18640 32036 18652
rect 32088 18640 32094 18692
rect 33594 18680 33600 18692
rect 33555 18652 33600 18680
rect 33594 18640 33600 18652
rect 33652 18640 33658 18692
rect 33796 18680 33824 18711
rect 33962 18708 33968 18760
rect 34020 18748 34026 18760
rect 34701 18751 34759 18757
rect 34701 18748 34713 18751
rect 34020 18720 34713 18748
rect 34020 18708 34026 18720
rect 34701 18717 34713 18720
rect 34747 18717 34759 18751
rect 34701 18711 34759 18717
rect 36078 18708 36084 18760
rect 36136 18708 36142 18760
rect 38764 18757 38792 18788
rect 40126 18776 40132 18788
rect 40184 18776 40190 18828
rect 43070 18776 43076 18828
rect 43128 18816 43134 18828
rect 47504 18825 47532 18924
rect 48593 18921 48605 18955
rect 48639 18952 48651 18955
rect 49694 18952 49700 18964
rect 48639 18924 49700 18952
rect 48639 18921 48651 18924
rect 48593 18915 48651 18921
rect 49694 18912 49700 18924
rect 49752 18912 49758 18964
rect 49786 18912 49792 18964
rect 49844 18952 49850 18964
rect 50341 18955 50399 18961
rect 50341 18952 50353 18955
rect 49844 18924 50353 18952
rect 49844 18912 49850 18924
rect 50341 18921 50353 18924
rect 50387 18952 50399 18955
rect 50522 18952 50528 18964
rect 50387 18924 50528 18952
rect 50387 18921 50399 18924
rect 50341 18915 50399 18921
rect 50522 18912 50528 18924
rect 50580 18912 50586 18964
rect 52181 18955 52239 18961
rect 52181 18921 52193 18955
rect 52227 18952 52239 18955
rect 52822 18952 52828 18964
rect 52227 18924 52828 18952
rect 52227 18921 52239 18924
rect 52181 18915 52239 18921
rect 52822 18912 52828 18924
rect 52880 18912 52886 18964
rect 53190 18952 53196 18964
rect 53151 18924 53196 18952
rect 53190 18912 53196 18924
rect 53248 18912 53254 18964
rect 49513 18887 49571 18893
rect 49513 18853 49525 18887
rect 49559 18884 49571 18887
rect 52638 18884 52644 18896
rect 49559 18856 52644 18884
rect 49559 18853 49571 18856
rect 49513 18847 49571 18853
rect 52638 18844 52644 18856
rect 52696 18844 52702 18896
rect 53101 18887 53159 18893
rect 53101 18853 53113 18887
rect 53147 18853 53159 18887
rect 53101 18847 53159 18853
rect 43257 18819 43315 18825
rect 43257 18816 43269 18819
rect 43128 18788 43269 18816
rect 43128 18776 43134 18788
rect 43257 18785 43269 18788
rect 43303 18785 43315 18819
rect 43257 18779 43315 18785
rect 47489 18819 47547 18825
rect 47489 18785 47501 18819
rect 47535 18785 47547 18819
rect 48406 18816 48412 18828
rect 48367 18788 48412 18816
rect 47489 18779 47547 18785
rect 48406 18776 48412 18788
rect 48464 18776 48470 18828
rect 52454 18816 52460 18828
rect 52104 18788 52460 18816
rect 37461 18751 37519 18757
rect 37461 18717 37473 18751
rect 37507 18717 37519 18751
rect 37461 18711 37519 18717
rect 38749 18751 38807 18757
rect 38749 18717 38761 18751
rect 38795 18717 38807 18751
rect 38749 18711 38807 18717
rect 34882 18680 34888 18692
rect 33796 18652 34888 18680
rect 34882 18640 34888 18652
rect 34940 18640 34946 18692
rect 34977 18683 35035 18689
rect 34977 18649 34989 18683
rect 35023 18649 35035 18683
rect 34977 18643 35035 18649
rect 24394 18612 24400 18624
rect 21284 18584 24400 18612
rect 24394 18572 24400 18584
rect 24452 18572 24458 18624
rect 26786 18612 26792 18624
rect 26747 18584 26792 18612
rect 26786 18572 26792 18584
rect 26844 18572 26850 18624
rect 29638 18572 29644 18624
rect 29696 18612 29702 18624
rect 34992 18612 35020 18643
rect 36262 18640 36268 18692
rect 36320 18680 36326 18692
rect 37476 18680 37504 18711
rect 39482 18708 39488 18760
rect 39540 18748 39546 18760
rect 39853 18751 39911 18757
rect 39853 18748 39865 18751
rect 39540 18720 39865 18748
rect 39540 18708 39546 18720
rect 39853 18717 39865 18720
rect 39899 18717 39911 18751
rect 39853 18711 39911 18717
rect 41230 18708 41236 18760
rect 41288 18708 41294 18760
rect 42426 18748 42432 18760
rect 42387 18720 42432 18748
rect 42426 18708 42432 18720
rect 42484 18708 42490 18760
rect 43530 18748 43536 18760
rect 43443 18720 43536 18748
rect 43530 18708 43536 18720
rect 43588 18748 43594 18760
rect 43990 18748 43996 18760
rect 43588 18720 43996 18748
rect 43588 18708 43594 18720
rect 43990 18708 43996 18720
rect 44048 18708 44054 18760
rect 44174 18748 44180 18760
rect 44135 18720 44180 18748
rect 44174 18708 44180 18720
rect 44232 18748 44238 18760
rect 46290 18748 46296 18760
rect 44232 18720 46296 18748
rect 44232 18708 44238 18720
rect 46290 18708 46296 18720
rect 46348 18708 46354 18760
rect 47670 18708 47676 18760
rect 47728 18748 47734 18760
rect 48317 18751 48375 18757
rect 48317 18748 48329 18751
rect 47728 18720 48329 18748
rect 47728 18708 47734 18720
rect 48317 18717 48329 18720
rect 48363 18748 48375 18751
rect 48682 18748 48688 18760
rect 48363 18720 48688 18748
rect 48363 18717 48375 18720
rect 48317 18711 48375 18717
rect 48682 18708 48688 18720
rect 48740 18708 48746 18760
rect 49329 18751 49387 18757
rect 49329 18717 49341 18751
rect 49375 18748 49387 18751
rect 50062 18748 50068 18760
rect 49375 18720 50068 18748
rect 49375 18717 49387 18720
rect 49329 18711 49387 18717
rect 50062 18708 50068 18720
rect 50120 18708 50126 18760
rect 52104 18757 52132 18788
rect 52454 18776 52460 18788
rect 52512 18816 52518 18828
rect 52914 18816 52920 18828
rect 52512 18788 52920 18816
rect 52512 18776 52518 18788
rect 52914 18776 52920 18788
rect 52972 18776 52978 18828
rect 53116 18816 53144 18847
rect 53190 18816 53196 18828
rect 53116 18788 53196 18816
rect 53190 18776 53196 18788
rect 53248 18776 53254 18828
rect 54754 18816 54760 18828
rect 54715 18788 54760 18816
rect 54754 18776 54760 18788
rect 54812 18776 54818 18828
rect 50157 18751 50215 18757
rect 50157 18717 50169 18751
rect 50203 18717 50215 18751
rect 50157 18711 50215 18717
rect 52089 18751 52147 18757
rect 52089 18717 52101 18751
rect 52135 18717 52147 18751
rect 52089 18711 52147 18717
rect 36320 18652 37504 18680
rect 38289 18683 38347 18689
rect 36320 18640 36326 18652
rect 38289 18649 38301 18683
rect 38335 18680 38347 18683
rect 42444 18680 42472 18708
rect 44453 18683 44511 18689
rect 38335 18652 39896 18680
rect 42444 18652 44404 18680
rect 38335 18649 38347 18652
rect 38289 18643 38347 18649
rect 29696 18584 35020 18612
rect 39868 18612 39896 18652
rect 41414 18612 41420 18624
rect 39868 18584 41420 18612
rect 29696 18572 29702 18584
rect 41414 18572 41420 18584
rect 41472 18572 41478 18624
rect 41598 18612 41604 18624
rect 41559 18584 41604 18612
rect 41598 18572 41604 18584
rect 41656 18572 41662 18624
rect 42521 18615 42579 18621
rect 42521 18581 42533 18615
rect 42567 18612 42579 18615
rect 42794 18612 42800 18624
rect 42567 18584 42800 18612
rect 42567 18581 42579 18584
rect 42521 18575 42579 18581
rect 42794 18572 42800 18584
rect 42852 18572 42858 18624
rect 44376 18612 44404 18652
rect 44453 18649 44465 18683
rect 44499 18680 44511 18683
rect 44634 18680 44640 18692
rect 44499 18652 44640 18680
rect 44499 18649 44511 18652
rect 44453 18643 44511 18649
rect 44634 18640 44640 18652
rect 44692 18640 44698 18692
rect 45189 18683 45247 18689
rect 45189 18649 45201 18683
rect 45235 18649 45247 18683
rect 45189 18643 45247 18649
rect 45833 18683 45891 18689
rect 45833 18649 45845 18683
rect 45879 18680 45891 18683
rect 45922 18680 45928 18692
rect 45879 18652 45928 18680
rect 45879 18649 45891 18652
rect 45833 18643 45891 18649
rect 45204 18612 45232 18643
rect 45922 18640 45928 18652
rect 45980 18640 45986 18692
rect 47394 18640 47400 18692
rect 47452 18680 47458 18692
rect 50172 18680 50200 18711
rect 52178 18708 52184 18760
rect 52236 18748 52242 18760
rect 52273 18751 52331 18757
rect 52273 18748 52285 18751
rect 52236 18720 52285 18748
rect 52236 18708 52242 18720
rect 52273 18717 52285 18720
rect 52319 18748 52331 18751
rect 54481 18751 54539 18757
rect 54481 18748 54493 18751
rect 52319 18720 54493 18748
rect 52319 18717 52331 18720
rect 52273 18711 52331 18717
rect 54481 18717 54493 18720
rect 54527 18717 54539 18751
rect 54481 18711 54539 18717
rect 57330 18708 57336 18760
rect 57388 18748 57394 18760
rect 57793 18751 57851 18757
rect 57793 18748 57805 18751
rect 57388 18720 57805 18748
rect 57388 18708 57394 18720
rect 57793 18717 57805 18720
rect 57839 18717 57851 18751
rect 57793 18711 57851 18717
rect 50798 18680 50804 18692
rect 47452 18652 50804 18680
rect 47452 18640 47458 18652
rect 50798 18640 50804 18652
rect 50856 18640 50862 18692
rect 52362 18640 52368 18692
rect 52420 18680 52426 18692
rect 52733 18683 52791 18689
rect 52733 18680 52745 18683
rect 52420 18652 52745 18680
rect 52420 18640 52426 18652
rect 52733 18649 52745 18652
rect 52779 18649 52791 18683
rect 52733 18643 52791 18649
rect 57422 18640 57428 18692
rect 57480 18680 57486 18692
rect 57609 18683 57667 18689
rect 57609 18680 57621 18683
rect 57480 18652 57621 18680
rect 57480 18640 57486 18652
rect 57609 18649 57621 18652
rect 57655 18649 57667 18683
rect 57609 18643 57667 18649
rect 44376 18584 45232 18612
rect 50893 18615 50951 18621
rect 50893 18581 50905 18615
rect 50939 18612 50951 18615
rect 51166 18612 51172 18624
rect 50939 18584 51172 18612
rect 50939 18581 50951 18584
rect 50893 18575 50951 18581
rect 51166 18572 51172 18584
rect 51224 18612 51230 18624
rect 51445 18615 51503 18621
rect 51445 18612 51457 18615
rect 51224 18584 51457 18612
rect 51224 18572 51230 18584
rect 51445 18581 51457 18584
rect 51491 18612 51503 18615
rect 54202 18612 54208 18624
rect 51491 18584 54208 18612
rect 51491 18581 51503 18584
rect 51445 18575 51503 18581
rect 54202 18572 54208 18584
rect 54260 18572 54266 18624
rect 1104 18522 58880 18544
rect 1104 18470 15398 18522
rect 15450 18470 15462 18522
rect 15514 18470 15526 18522
rect 15578 18470 15590 18522
rect 15642 18470 15654 18522
rect 15706 18470 29846 18522
rect 29898 18470 29910 18522
rect 29962 18470 29974 18522
rect 30026 18470 30038 18522
rect 30090 18470 30102 18522
rect 30154 18470 44294 18522
rect 44346 18470 44358 18522
rect 44410 18470 44422 18522
rect 44474 18470 44486 18522
rect 44538 18470 44550 18522
rect 44602 18470 58880 18522
rect 1104 18448 58880 18470
rect 4249 18411 4307 18417
rect 4249 18377 4261 18411
rect 4295 18408 4307 18411
rect 4338 18408 4344 18420
rect 4295 18380 4344 18408
rect 4295 18377 4307 18380
rect 4249 18371 4307 18377
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 5074 18408 5080 18420
rect 5035 18380 5080 18408
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 5721 18411 5779 18417
rect 5721 18377 5733 18411
rect 5767 18408 5779 18411
rect 6270 18408 6276 18420
rect 5767 18380 6276 18408
rect 5767 18377 5779 18380
rect 5721 18371 5779 18377
rect 6270 18368 6276 18380
rect 6328 18368 6334 18420
rect 7006 18368 7012 18420
rect 7064 18368 7070 18420
rect 10226 18368 10232 18420
rect 10284 18408 10290 18420
rect 11238 18408 11244 18420
rect 10284 18380 11244 18408
rect 10284 18368 10290 18380
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 14642 18408 14648 18420
rect 14603 18380 14648 18408
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 15565 18411 15623 18417
rect 15565 18377 15577 18411
rect 15611 18408 15623 18411
rect 16482 18408 16488 18420
rect 15611 18380 16488 18408
rect 15611 18377 15623 18380
rect 15565 18371 15623 18377
rect 16482 18368 16488 18380
rect 16540 18408 16546 18420
rect 19518 18408 19524 18420
rect 16540 18380 19524 18408
rect 16540 18368 16546 18380
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 21174 18408 21180 18420
rect 21135 18380 21180 18408
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 22094 18408 22100 18420
rect 22066 18368 22100 18408
rect 22152 18368 22158 18420
rect 24854 18408 24860 18420
rect 23952 18380 24860 18408
rect 4706 18300 4712 18352
rect 4764 18340 4770 18352
rect 4764 18312 6960 18340
rect 4764 18300 4770 18312
rect 2130 18272 2136 18284
rect 2091 18244 2136 18272
rect 2130 18232 2136 18244
rect 2188 18232 2194 18284
rect 3881 18275 3939 18281
rect 3881 18241 3893 18275
rect 3927 18272 3939 18275
rect 4062 18272 4068 18284
rect 3927 18244 4068 18272
rect 3927 18241 3939 18244
rect 3881 18235 3939 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 5169 18275 5227 18281
rect 5169 18241 5181 18275
rect 5215 18241 5227 18275
rect 5626 18272 5632 18284
rect 5587 18244 5632 18272
rect 5169 18235 5227 18241
rect 2222 18204 2228 18216
rect 2183 18176 2228 18204
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 3786 18204 3792 18216
rect 2915 18176 3792 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 3970 18204 3976 18216
rect 3931 18176 3976 18204
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 5184 18204 5212 18235
rect 5626 18232 5632 18244
rect 5684 18232 5690 18284
rect 5902 18232 5908 18284
rect 5960 18272 5966 18284
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 5960 18244 6377 18272
rect 5960 18232 5966 18244
rect 6365 18241 6377 18244
rect 6411 18272 6423 18275
rect 6411 18244 6868 18272
rect 6411 18241 6423 18244
rect 6365 18235 6423 18241
rect 6270 18204 6276 18216
rect 5184 18176 6276 18204
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 6454 18068 6460 18080
rect 6415 18040 6460 18068
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 6840 18068 6868 18244
rect 6932 18204 6960 18312
rect 7024 18281 7052 18368
rect 7282 18300 7288 18352
rect 7340 18340 7346 18352
rect 10965 18343 11023 18349
rect 7340 18312 7774 18340
rect 7340 18300 7346 18312
rect 10965 18309 10977 18343
rect 11011 18340 11023 18343
rect 13078 18340 13084 18352
rect 11011 18312 13084 18340
rect 11011 18309 11023 18312
rect 10965 18303 11023 18309
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 13262 18300 13268 18352
rect 13320 18340 13326 18352
rect 18414 18340 18420 18352
rect 13320 18312 16712 18340
rect 18170 18312 18420 18340
rect 13320 18300 13326 18312
rect 6998 18275 7056 18281
rect 6998 18241 7010 18275
rect 7044 18241 7056 18275
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 6998 18235 7056 18241
rect 9692 18244 11529 18272
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6932 18176 7297 18204
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 9692 18145 9720 18244
rect 11517 18241 11529 18244
rect 11563 18272 11575 18275
rect 11698 18272 11704 18284
rect 11563 18244 11704 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 12253 18275 12311 18281
rect 12253 18241 12265 18275
rect 12299 18241 12311 18275
rect 13170 18272 13176 18284
rect 13131 18244 13176 18272
rect 12253 18235 12311 18241
rect 11330 18164 11336 18216
rect 11388 18204 11394 18216
rect 12268 18204 12296 18235
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 14734 18272 14740 18284
rect 14695 18244 14740 18272
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 16684 18281 16712 18312
rect 18414 18300 18420 18312
rect 18472 18300 18478 18352
rect 18690 18300 18696 18352
rect 18748 18340 18754 18352
rect 22066 18340 22094 18368
rect 23952 18349 23980 18380
rect 24854 18368 24860 18380
rect 24912 18368 24918 18420
rect 25038 18368 25044 18420
rect 25096 18408 25102 18420
rect 27249 18411 27307 18417
rect 27249 18408 27261 18411
rect 25096 18380 27261 18408
rect 25096 18368 25102 18380
rect 27249 18377 27261 18380
rect 27295 18408 27307 18411
rect 28077 18411 28135 18417
rect 28077 18408 28089 18411
rect 27295 18380 28089 18408
rect 27295 18377 27307 18380
rect 27249 18371 27307 18377
rect 28077 18377 28089 18380
rect 28123 18377 28135 18411
rect 28077 18371 28135 18377
rect 29549 18411 29607 18417
rect 29549 18377 29561 18411
rect 29595 18408 29607 18411
rect 29638 18408 29644 18420
rect 29595 18380 29644 18408
rect 29595 18377 29607 18380
rect 29549 18371 29607 18377
rect 29638 18368 29644 18380
rect 29696 18368 29702 18420
rect 30190 18368 30196 18420
rect 30248 18408 30254 18420
rect 33962 18408 33968 18420
rect 30248 18380 33968 18408
rect 30248 18368 30254 18380
rect 33962 18368 33968 18380
rect 34020 18368 34026 18420
rect 34882 18368 34888 18420
rect 34940 18408 34946 18420
rect 34940 18380 35388 18408
rect 34940 18368 34946 18380
rect 18748 18312 22094 18340
rect 23937 18343 23995 18349
rect 18748 18300 18754 18312
rect 23937 18309 23949 18343
rect 23983 18309 23995 18343
rect 24946 18340 24952 18352
rect 23937 18303 23995 18309
rect 24044 18312 24952 18340
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18241 16727 18275
rect 18966 18272 18972 18284
rect 18927 18244 18972 18272
rect 16669 18235 16727 18241
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19116 18244 19380 18272
rect 19116 18232 19122 18244
rect 11388 18176 12296 18204
rect 16945 18207 17003 18213
rect 11388 18164 11394 18176
rect 16945 18173 16957 18207
rect 16991 18204 17003 18207
rect 18690 18204 18696 18216
rect 16991 18176 18696 18204
rect 16991 18173 17003 18176
rect 16945 18167 17003 18173
rect 18690 18164 18696 18176
rect 18748 18164 18754 18216
rect 19352 18204 19380 18244
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 22189 18275 22247 18281
rect 22189 18272 22201 18275
rect 22152 18244 22201 18272
rect 22152 18232 22158 18244
rect 22189 18241 22201 18244
rect 22235 18272 22247 18275
rect 24044 18272 24072 18312
rect 24946 18300 24952 18312
rect 25004 18300 25010 18352
rect 25682 18300 25688 18352
rect 25740 18300 25746 18352
rect 26050 18300 26056 18352
rect 26108 18340 26114 18352
rect 30650 18340 30656 18352
rect 26108 18312 30656 18340
rect 26108 18300 26114 18312
rect 30650 18300 30656 18312
rect 30708 18300 30714 18352
rect 30837 18343 30895 18349
rect 30837 18309 30849 18343
rect 30883 18340 30895 18343
rect 31938 18340 31944 18352
rect 30883 18312 31944 18340
rect 30883 18309 30895 18312
rect 30837 18303 30895 18309
rect 31938 18300 31944 18312
rect 31996 18300 32002 18352
rect 33870 18340 33876 18352
rect 32324 18312 33876 18340
rect 22235 18244 24072 18272
rect 27157 18275 27215 18281
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 27157 18241 27169 18275
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18272 27399 18275
rect 27430 18272 27436 18284
rect 27387 18244 27436 18272
rect 27387 18241 27399 18244
rect 27341 18235 27399 18241
rect 24397 18207 24455 18213
rect 24397 18204 24409 18207
rect 19352 18176 24409 18204
rect 24397 18173 24409 18176
rect 24443 18173 24455 18207
rect 24670 18204 24676 18216
rect 24631 18176 24676 18204
rect 24397 18167 24455 18173
rect 24670 18164 24676 18176
rect 24728 18164 24734 18216
rect 25222 18164 25228 18216
rect 25280 18204 25286 18216
rect 26142 18204 26148 18216
rect 25280 18176 26148 18204
rect 25280 18164 25286 18176
rect 26142 18164 26148 18176
rect 26200 18164 26206 18216
rect 27172 18204 27200 18235
rect 27430 18232 27436 18244
rect 27488 18232 27494 18284
rect 28166 18272 28172 18284
rect 27724 18244 28172 18272
rect 27724 18216 27752 18244
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 29181 18275 29239 18281
rect 29181 18272 29193 18275
rect 28460 18244 29193 18272
rect 27706 18204 27712 18216
rect 27172 18176 27712 18204
rect 27706 18164 27712 18176
rect 27764 18164 27770 18216
rect 27985 18207 28043 18213
rect 27985 18173 27997 18207
rect 28031 18204 28043 18207
rect 28074 18204 28080 18216
rect 28031 18176 28080 18204
rect 28031 18173 28043 18176
rect 27985 18167 28043 18173
rect 28074 18164 28080 18176
rect 28132 18164 28138 18216
rect 9677 18139 9735 18145
rect 9677 18105 9689 18139
rect 9723 18105 9735 18139
rect 9677 18099 9735 18105
rect 11974 18096 11980 18148
rect 12032 18136 12038 18148
rect 16022 18136 16028 18148
rect 12032 18108 16028 18136
rect 12032 18096 12038 18108
rect 16022 18096 16028 18108
rect 16080 18096 16086 18148
rect 18417 18139 18475 18145
rect 18417 18105 18429 18139
rect 18463 18136 18475 18139
rect 21818 18136 21824 18148
rect 18463 18108 21824 18136
rect 18463 18105 18475 18108
rect 18417 18099 18475 18105
rect 21818 18096 21824 18108
rect 21876 18096 21882 18148
rect 26234 18096 26240 18148
rect 26292 18136 26298 18148
rect 28460 18136 28488 18244
rect 29181 18241 29193 18244
rect 29227 18272 29239 18275
rect 30466 18272 30472 18284
rect 29227 18244 30472 18272
rect 29227 18241 29239 18244
rect 29181 18235 29239 18241
rect 30466 18232 30472 18244
rect 30524 18232 30530 18284
rect 30926 18272 30932 18284
rect 30839 18244 30932 18272
rect 30926 18232 30932 18244
rect 30984 18272 30990 18284
rect 31110 18272 31116 18284
rect 30984 18244 31116 18272
rect 30984 18232 30990 18244
rect 31110 18232 31116 18244
rect 31168 18232 31174 18284
rect 31202 18232 31208 18284
rect 31260 18272 31266 18284
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 31260 18244 31493 18272
rect 31260 18232 31266 18244
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 31481 18235 31539 18241
rect 31573 18275 31631 18281
rect 31573 18241 31585 18275
rect 31619 18272 31631 18275
rect 32324 18272 32352 18312
rect 33870 18300 33876 18312
rect 33928 18300 33934 18352
rect 35158 18340 35164 18352
rect 34440 18312 35164 18340
rect 32582 18272 32588 18284
rect 31619 18244 32352 18272
rect 32543 18244 32588 18272
rect 31619 18241 31631 18244
rect 31573 18235 31631 18241
rect 32582 18232 32588 18244
rect 32640 18232 32646 18284
rect 33134 18232 33140 18284
rect 33192 18272 33198 18284
rect 34440 18281 34468 18312
rect 35158 18300 35164 18312
rect 35216 18300 35222 18352
rect 35360 18340 35388 18380
rect 35434 18368 35440 18420
rect 35492 18408 35498 18420
rect 41046 18408 41052 18420
rect 35492 18380 40448 18408
rect 41007 18380 41052 18408
rect 35492 18368 35498 18380
rect 36538 18340 36544 18352
rect 35360 18312 36544 18340
rect 36538 18300 36544 18312
rect 36596 18300 36602 18352
rect 38378 18300 38384 18352
rect 38436 18340 38442 18352
rect 40313 18343 40371 18349
rect 40313 18340 40325 18343
rect 38436 18312 40325 18340
rect 38436 18300 38442 18312
rect 40313 18309 40325 18312
rect 40359 18309 40371 18343
rect 40420 18340 40448 18380
rect 41046 18368 41052 18380
rect 41104 18368 41110 18420
rect 48774 18408 48780 18420
rect 41386 18380 48780 18408
rect 41386 18340 41414 18380
rect 48774 18368 48780 18380
rect 48832 18368 48838 18420
rect 49602 18408 49608 18420
rect 49252 18380 49608 18408
rect 40420 18312 41414 18340
rect 40313 18303 40371 18309
rect 42058 18300 42064 18352
rect 42116 18340 42122 18352
rect 42116 18312 42472 18340
rect 42116 18300 42122 18312
rect 33229 18275 33287 18281
rect 33229 18272 33241 18275
rect 33192 18244 33241 18272
rect 33192 18232 33198 18244
rect 33229 18241 33241 18244
rect 33275 18272 33287 18275
rect 34425 18275 34483 18281
rect 33275 18244 34376 18272
rect 33275 18241 33287 18244
rect 33229 18235 33287 18241
rect 29270 18204 29276 18216
rect 28552 18176 29276 18204
rect 28552 18145 28580 18176
rect 29270 18164 29276 18176
rect 29328 18164 29334 18216
rect 32677 18207 32735 18213
rect 32677 18173 32689 18207
rect 32723 18204 32735 18207
rect 34238 18204 34244 18216
rect 32723 18176 34244 18204
rect 32723 18173 32735 18176
rect 32677 18167 32735 18173
rect 34238 18164 34244 18176
rect 34296 18164 34302 18216
rect 26292 18108 28488 18136
rect 28537 18139 28595 18145
rect 26292 18096 26298 18108
rect 28537 18105 28549 18139
rect 28583 18105 28595 18139
rect 34348 18136 34376 18244
rect 34425 18241 34437 18275
rect 34471 18241 34483 18275
rect 38470 18272 38476 18284
rect 34425 18235 34483 18241
rect 37844 18244 38476 18272
rect 34606 18204 34612 18216
rect 34567 18176 34612 18204
rect 34606 18164 34612 18176
rect 34664 18164 34670 18216
rect 34790 18164 34796 18216
rect 34848 18204 34854 18216
rect 34885 18207 34943 18213
rect 34885 18204 34897 18207
rect 34848 18176 34897 18204
rect 34848 18164 34854 18176
rect 34885 18173 34897 18176
rect 34931 18173 34943 18207
rect 34885 18167 34943 18173
rect 36446 18164 36452 18216
rect 36504 18204 36510 18216
rect 37844 18213 37872 18244
rect 38470 18232 38476 18244
rect 38528 18232 38534 18284
rect 40862 18232 40868 18284
rect 40920 18272 40926 18284
rect 40957 18275 41015 18281
rect 40957 18272 40969 18275
rect 40920 18244 40969 18272
rect 40920 18232 40926 18244
rect 40957 18241 40969 18244
rect 41003 18241 41015 18275
rect 40957 18235 41015 18241
rect 41601 18275 41659 18281
rect 41601 18241 41613 18275
rect 41647 18272 41659 18275
rect 41690 18272 41696 18284
rect 41647 18244 41696 18272
rect 41647 18241 41659 18244
rect 41601 18235 41659 18241
rect 41690 18232 41696 18244
rect 41748 18232 41754 18284
rect 42444 18281 42472 18312
rect 42518 18300 42524 18352
rect 42576 18340 42582 18352
rect 42576 18312 44496 18340
rect 42576 18300 42582 18312
rect 42429 18275 42487 18281
rect 42429 18241 42441 18275
rect 42475 18241 42487 18275
rect 42429 18235 42487 18241
rect 42610 18232 42616 18284
rect 42668 18272 42674 18284
rect 42705 18275 42763 18281
rect 42705 18272 42717 18275
rect 42668 18244 42717 18272
rect 42668 18232 42674 18244
rect 42705 18241 42717 18244
rect 42751 18241 42763 18275
rect 43346 18272 43352 18284
rect 43307 18244 43352 18272
rect 42705 18235 42763 18241
rect 43346 18232 43352 18244
rect 43404 18232 43410 18284
rect 44468 18281 44496 18312
rect 44634 18300 44640 18352
rect 44692 18340 44698 18352
rect 45554 18340 45560 18352
rect 44692 18312 45560 18340
rect 44692 18300 44698 18312
rect 45554 18300 45560 18312
rect 45612 18300 45618 18352
rect 45830 18300 45836 18352
rect 45888 18340 45894 18352
rect 48041 18343 48099 18349
rect 48041 18340 48053 18343
rect 45888 18312 48053 18340
rect 45888 18300 45894 18312
rect 48041 18309 48053 18312
rect 48087 18309 48099 18343
rect 48041 18303 48099 18309
rect 48225 18343 48283 18349
rect 48225 18309 48237 18343
rect 48271 18340 48283 18343
rect 49252 18340 49280 18380
rect 49602 18368 49608 18380
rect 49660 18408 49666 18420
rect 49660 18380 50200 18408
rect 49660 18368 49666 18380
rect 50172 18340 50200 18380
rect 50246 18340 50252 18352
rect 48271 18312 49280 18340
rect 50094 18312 50252 18340
rect 48271 18309 48283 18312
rect 48225 18303 48283 18309
rect 50246 18300 50252 18312
rect 50304 18300 50310 18352
rect 52730 18300 52736 18352
rect 52788 18340 52794 18352
rect 52788 18312 53052 18340
rect 52788 18300 52794 18312
rect 44453 18275 44511 18281
rect 44453 18241 44465 18275
rect 44499 18241 44511 18275
rect 44453 18235 44511 18241
rect 50798 18232 50804 18284
rect 50856 18272 50862 18284
rect 50856 18244 50901 18272
rect 50856 18232 50862 18244
rect 51074 18232 51080 18284
rect 51132 18272 51138 18284
rect 51261 18275 51319 18281
rect 51261 18272 51273 18275
rect 51132 18244 51273 18272
rect 51132 18232 51138 18244
rect 51261 18241 51273 18244
rect 51307 18241 51319 18275
rect 51261 18235 51319 18241
rect 51445 18275 51503 18281
rect 51445 18241 51457 18275
rect 51491 18241 51503 18275
rect 51994 18272 52000 18284
rect 51955 18244 52000 18272
rect 51445 18235 51503 18241
rect 37829 18207 37887 18213
rect 37829 18204 37841 18207
rect 36504 18176 37841 18204
rect 36504 18164 36510 18176
rect 37829 18173 37841 18176
rect 37875 18173 37887 18207
rect 38102 18204 38108 18216
rect 38063 18176 38108 18204
rect 37829 18167 37887 18173
rect 38102 18164 38108 18176
rect 38160 18164 38166 18216
rect 40037 18207 40095 18213
rect 40037 18173 40049 18207
rect 40083 18173 40095 18207
rect 40037 18167 40095 18173
rect 40497 18207 40555 18213
rect 40497 18173 40509 18207
rect 40543 18173 40555 18207
rect 40497 18167 40555 18173
rect 34698 18136 34704 18148
rect 34348 18108 34704 18136
rect 28537 18099 28595 18105
rect 34698 18096 34704 18108
rect 34756 18096 34762 18148
rect 8570 18068 8576 18080
rect 6840 18040 8576 18068
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 8757 18071 8815 18077
rect 8757 18037 8769 18071
rect 8803 18068 8815 18071
rect 9214 18068 9220 18080
rect 8803 18040 9220 18068
rect 8803 18037 8815 18040
rect 8757 18031 8815 18037
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 11606 18068 11612 18080
rect 11567 18040 11612 18068
rect 11606 18028 11612 18040
rect 11664 18028 11670 18080
rect 14090 18068 14096 18080
rect 14051 18040 14096 18068
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 20254 18068 20260 18080
rect 20215 18040 20260 18068
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 21174 18028 21180 18080
rect 21232 18068 21238 18080
rect 22462 18068 22468 18080
rect 21232 18040 22468 18068
rect 21232 18028 21238 18040
rect 22462 18028 22468 18040
rect 22520 18028 22526 18080
rect 33226 18068 33232 18080
rect 33187 18040 33232 18068
rect 33226 18028 33232 18040
rect 33284 18028 33290 18080
rect 33962 18068 33968 18080
rect 33923 18040 33968 18068
rect 33962 18028 33968 18040
rect 34020 18028 34026 18080
rect 34238 18028 34244 18080
rect 34296 18068 34302 18080
rect 39482 18068 39488 18080
rect 34296 18040 39488 18068
rect 34296 18028 34302 18040
rect 39482 18028 39488 18040
rect 39540 18028 39546 18080
rect 40052 18068 40080 18167
rect 40512 18136 40540 18167
rect 41414 18164 41420 18216
rect 41472 18204 41478 18216
rect 42334 18204 42340 18216
rect 41472 18176 42340 18204
rect 41472 18164 41478 18176
rect 42334 18164 42340 18176
rect 42392 18164 42398 18216
rect 44545 18207 44603 18213
rect 44545 18173 44557 18207
rect 44591 18173 44603 18207
rect 45922 18204 45928 18216
rect 45883 18176 45928 18204
rect 44545 18167 44603 18173
rect 42426 18136 42432 18148
rect 40512 18108 42432 18136
rect 42426 18096 42432 18108
rect 42484 18096 42490 18148
rect 43806 18096 43812 18148
rect 43864 18136 43870 18148
rect 44085 18139 44143 18145
rect 44085 18136 44097 18139
rect 43864 18108 44097 18136
rect 43864 18096 43870 18108
rect 44085 18105 44097 18108
rect 44131 18105 44143 18139
rect 44560 18136 44588 18167
rect 45922 18164 45928 18176
rect 45980 18164 45986 18216
rect 46842 18204 46848 18216
rect 46803 18176 46848 18204
rect 46842 18164 46848 18176
rect 46900 18164 46906 18216
rect 47026 18204 47032 18216
rect 46987 18176 47032 18204
rect 47026 18164 47032 18176
rect 47084 18164 47090 18216
rect 50062 18204 50068 18216
rect 48700 18176 50068 18204
rect 46750 18136 46756 18148
rect 44560 18108 46756 18136
rect 44085 18099 44143 18105
rect 46750 18096 46756 18108
rect 46808 18096 46814 18148
rect 46860 18136 46888 18164
rect 48590 18136 48596 18148
rect 46860 18108 48596 18136
rect 48590 18096 48596 18108
rect 48648 18096 48654 18148
rect 41414 18068 41420 18080
rect 40052 18040 41420 18068
rect 41414 18028 41420 18040
rect 41472 18028 41478 18080
rect 41785 18071 41843 18077
rect 41785 18037 41797 18071
rect 41831 18068 41843 18071
rect 42978 18068 42984 18080
rect 41831 18040 42984 18068
rect 41831 18037 41843 18040
rect 41785 18031 41843 18037
rect 42978 18028 42984 18040
rect 43036 18028 43042 18080
rect 43625 18071 43683 18077
rect 43625 18037 43637 18071
rect 43671 18068 43683 18071
rect 43990 18068 43996 18080
rect 43671 18040 43996 18068
rect 43671 18037 43683 18040
rect 43625 18031 43683 18037
rect 43990 18028 43996 18040
rect 44048 18068 44054 18080
rect 48700 18068 48728 18176
rect 50062 18164 50068 18176
rect 50120 18164 50126 18216
rect 50522 18204 50528 18216
rect 50483 18176 50528 18204
rect 50522 18164 50528 18176
rect 50580 18164 50586 18216
rect 51460 18204 51488 18235
rect 51994 18232 52000 18244
rect 52052 18232 52058 18284
rect 52178 18272 52184 18284
rect 52139 18244 52184 18272
rect 52178 18232 52184 18244
rect 52236 18272 52242 18284
rect 52822 18272 52828 18284
rect 52236 18244 52828 18272
rect 52236 18232 52242 18244
rect 52822 18232 52828 18244
rect 52880 18232 52886 18284
rect 53024 18281 53052 18312
rect 53009 18275 53067 18281
rect 53009 18241 53021 18275
rect 53055 18272 53067 18275
rect 53282 18272 53288 18284
rect 53055 18244 53288 18272
rect 53055 18241 53067 18244
rect 53009 18235 53067 18241
rect 53282 18232 53288 18244
rect 53340 18272 53346 18284
rect 54573 18275 54631 18281
rect 54573 18272 54585 18275
rect 53340 18244 54585 18272
rect 53340 18232 53346 18244
rect 54573 18241 54585 18244
rect 54619 18241 54631 18275
rect 54573 18235 54631 18241
rect 56321 18275 56379 18281
rect 56321 18241 56333 18275
rect 56367 18272 56379 18275
rect 56410 18272 56416 18284
rect 56367 18244 56416 18272
rect 56367 18241 56379 18244
rect 56321 18235 56379 18241
rect 56410 18232 56416 18244
rect 56468 18232 56474 18284
rect 57882 18272 57888 18284
rect 57843 18244 57888 18272
rect 57882 18232 57888 18244
rect 57940 18232 57946 18284
rect 52733 18207 52791 18213
rect 52733 18204 52745 18207
rect 51460 18176 52745 18204
rect 52733 18173 52745 18176
rect 52779 18173 52791 18207
rect 52733 18167 52791 18173
rect 52917 18207 52975 18213
rect 52917 18173 52929 18207
rect 52963 18204 52975 18207
rect 53101 18207 53159 18213
rect 52963 18176 53052 18204
rect 52963 18173 52975 18176
rect 52917 18167 52975 18173
rect 53024 18148 53052 18176
rect 53101 18173 53113 18207
rect 53147 18173 53159 18207
rect 53101 18167 53159 18173
rect 53006 18096 53012 18148
rect 53064 18096 53070 18148
rect 53116 18136 53144 18167
rect 53190 18164 53196 18216
rect 53248 18204 53254 18216
rect 53248 18176 53293 18204
rect 53248 18164 53254 18176
rect 54110 18164 54116 18216
rect 54168 18204 54174 18216
rect 54297 18207 54355 18213
rect 54297 18204 54309 18207
rect 54168 18176 54309 18204
rect 54168 18164 54174 18176
rect 54297 18173 54309 18176
rect 54343 18173 54355 18207
rect 56226 18204 56232 18216
rect 56187 18176 56232 18204
rect 54297 18167 54355 18173
rect 56226 18164 56232 18176
rect 56284 18164 56290 18216
rect 53466 18136 53472 18148
rect 53116 18108 53472 18136
rect 53466 18096 53472 18108
rect 53524 18096 53530 18148
rect 56686 18136 56692 18148
rect 56647 18108 56692 18136
rect 56686 18096 56692 18108
rect 56744 18096 56750 18148
rect 49050 18068 49056 18080
rect 44048 18040 48728 18068
rect 49011 18040 49056 18068
rect 44048 18028 44054 18040
rect 49050 18028 49056 18040
rect 49108 18028 49114 18080
rect 50430 18028 50436 18080
rect 50488 18068 50494 18080
rect 51353 18071 51411 18077
rect 51353 18068 51365 18071
rect 50488 18040 51365 18068
rect 50488 18028 50494 18040
rect 51353 18037 51365 18040
rect 51399 18037 51411 18071
rect 51353 18031 51411 18037
rect 52089 18071 52147 18077
rect 52089 18037 52101 18071
rect 52135 18068 52147 18071
rect 53558 18068 53564 18080
rect 52135 18040 53564 18068
rect 52135 18037 52147 18040
rect 52089 18031 52147 18037
rect 53558 18028 53564 18040
rect 53616 18028 53622 18080
rect 53834 18068 53840 18080
rect 53747 18040 53840 18068
rect 53834 18028 53840 18040
rect 53892 18068 53898 18080
rect 55950 18068 55956 18080
rect 53892 18040 55956 18068
rect 53892 18028 53898 18040
rect 55950 18028 55956 18040
rect 56008 18028 56014 18080
rect 57790 18028 57796 18080
rect 57848 18068 57854 18080
rect 58069 18071 58127 18077
rect 58069 18068 58081 18071
rect 57848 18040 58081 18068
rect 57848 18028 57854 18040
rect 58069 18037 58081 18040
rect 58115 18037 58127 18071
rect 58069 18031 58127 18037
rect 1104 17978 58880 18000
rect 1104 17926 8174 17978
rect 8226 17926 8238 17978
rect 8290 17926 8302 17978
rect 8354 17926 8366 17978
rect 8418 17926 8430 17978
rect 8482 17926 22622 17978
rect 22674 17926 22686 17978
rect 22738 17926 22750 17978
rect 22802 17926 22814 17978
rect 22866 17926 22878 17978
rect 22930 17926 37070 17978
rect 37122 17926 37134 17978
rect 37186 17926 37198 17978
rect 37250 17926 37262 17978
rect 37314 17926 37326 17978
rect 37378 17926 51518 17978
rect 51570 17926 51582 17978
rect 51634 17926 51646 17978
rect 51698 17926 51710 17978
rect 51762 17926 51774 17978
rect 51826 17926 58880 17978
rect 1104 17904 58880 17926
rect 2130 17824 2136 17876
rect 2188 17864 2194 17876
rect 3053 17867 3111 17873
rect 3053 17864 3065 17867
rect 2188 17836 3065 17864
rect 2188 17824 2194 17836
rect 3053 17833 3065 17836
rect 3099 17833 3111 17867
rect 3053 17827 3111 17833
rect 9033 17867 9091 17873
rect 9033 17833 9045 17867
rect 9079 17864 9091 17867
rect 11054 17864 11060 17876
rect 9079 17836 11060 17864
rect 9079 17833 9091 17836
rect 9033 17827 9091 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 11333 17867 11391 17873
rect 11333 17833 11345 17867
rect 11379 17864 11391 17867
rect 11422 17864 11428 17876
rect 11379 17836 11428 17864
rect 11379 17833 11391 17836
rect 11333 17827 11391 17833
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 16206 17864 16212 17876
rect 15344 17836 16212 17864
rect 15344 17824 15350 17836
rect 16206 17824 16212 17836
rect 16264 17864 16270 17876
rect 20254 17864 20260 17876
rect 16264 17836 20260 17864
rect 16264 17824 16270 17836
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 22833 17867 22891 17873
rect 22833 17833 22845 17867
rect 22879 17864 22891 17867
rect 22922 17864 22928 17876
rect 22879 17836 22928 17864
rect 22879 17833 22891 17836
rect 22833 17827 22891 17833
rect 22922 17824 22928 17836
rect 22980 17824 22986 17876
rect 23014 17824 23020 17876
rect 23072 17864 23078 17876
rect 23566 17864 23572 17876
rect 23072 17836 23572 17864
rect 23072 17824 23078 17836
rect 23566 17824 23572 17836
rect 23624 17824 23630 17876
rect 24946 17824 24952 17876
rect 25004 17864 25010 17876
rect 26237 17867 26295 17873
rect 26237 17864 26249 17867
rect 25004 17836 26249 17864
rect 25004 17824 25010 17836
rect 26237 17833 26249 17836
rect 26283 17833 26295 17867
rect 26237 17827 26295 17833
rect 36814 17824 36820 17876
rect 36872 17864 36878 17876
rect 38286 17864 38292 17876
rect 36872 17836 38292 17864
rect 36872 17824 36878 17836
rect 38286 17824 38292 17836
rect 38344 17824 38350 17876
rect 41414 17824 41420 17876
rect 41472 17864 41478 17876
rect 41601 17867 41659 17873
rect 41601 17864 41613 17867
rect 41472 17836 41613 17864
rect 41472 17824 41478 17836
rect 41601 17833 41613 17836
rect 41647 17864 41659 17867
rect 41874 17864 41880 17876
rect 41647 17836 41880 17864
rect 41647 17833 41659 17836
rect 41601 17827 41659 17833
rect 41874 17824 41880 17836
rect 41932 17824 41938 17876
rect 42383 17867 42441 17873
rect 42383 17833 42395 17867
rect 42429 17864 42441 17867
rect 42518 17864 42524 17876
rect 42429 17836 42524 17864
rect 42429 17833 42441 17836
rect 42383 17827 42441 17833
rect 42518 17824 42524 17836
rect 42576 17824 42582 17876
rect 50522 17824 50528 17876
rect 50580 17864 50586 17876
rect 50617 17867 50675 17873
rect 50617 17864 50629 17867
rect 50580 17836 50629 17864
rect 50580 17824 50586 17836
rect 50617 17833 50629 17836
rect 50663 17833 50675 17867
rect 52178 17864 52184 17876
rect 50617 17827 50675 17833
rect 51046 17836 52184 17864
rect 4246 17796 4252 17808
rect 3252 17768 4252 17796
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17728 2283 17731
rect 2866 17728 2872 17740
rect 2271 17700 2872 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 3050 17660 3056 17672
rect 2179 17632 3056 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 3252 17669 3280 17768
rect 4246 17756 4252 17768
rect 4304 17756 4310 17808
rect 11514 17796 11520 17808
rect 10888 17768 11520 17796
rect 5166 17688 5172 17740
rect 5224 17728 5230 17740
rect 6825 17731 6883 17737
rect 6825 17728 6837 17731
rect 5224 17700 6837 17728
rect 5224 17688 5230 17700
rect 6825 17697 6837 17700
rect 6871 17697 6883 17731
rect 10888 17728 10916 17768
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 11882 17756 11888 17808
rect 11940 17796 11946 17808
rect 18598 17796 18604 17808
rect 11940 17768 14872 17796
rect 18559 17768 18604 17796
rect 11940 17756 11946 17768
rect 14844 17737 14872 17768
rect 18598 17756 18604 17768
rect 18656 17756 18662 17808
rect 18690 17756 18696 17808
rect 18748 17796 18754 17808
rect 19797 17799 19855 17805
rect 19797 17796 19809 17799
rect 18748 17768 19809 17796
rect 18748 17756 18754 17768
rect 19797 17765 19809 17768
rect 19843 17765 19855 17799
rect 23477 17799 23535 17805
rect 19797 17759 19855 17765
rect 19904 17768 22876 17796
rect 14185 17731 14243 17737
rect 14185 17728 14197 17731
rect 6825 17691 6883 17697
rect 9140 17700 10916 17728
rect 11624 17700 14197 17728
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17629 3295 17663
rect 4798 17660 4804 17672
rect 4759 17632 4804 17660
rect 3237 17623 3295 17629
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 5077 17663 5135 17669
rect 5077 17629 5089 17663
rect 5123 17660 5135 17663
rect 5626 17660 5632 17672
rect 5123 17632 5632 17660
rect 5123 17629 5135 17632
rect 5077 17623 5135 17629
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 9140 17669 9168 17700
rect 6549 17663 6607 17669
rect 6549 17629 6561 17663
rect 6595 17629 6607 17663
rect 6549 17623 6607 17629
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17629 9183 17663
rect 9582 17660 9588 17672
rect 9543 17632 9588 17660
rect 9125 17623 9183 17629
rect 5718 17592 5724 17604
rect 5679 17564 5724 17592
rect 5718 17552 5724 17564
rect 5776 17552 5782 17604
rect 6564 17592 6592 17623
rect 9582 17620 9588 17632
rect 9640 17620 9646 17672
rect 11624 17660 11652 17700
rect 14185 17697 14197 17700
rect 14231 17697 14243 17731
rect 14185 17691 14243 17697
rect 14829 17731 14887 17737
rect 14829 17697 14841 17731
rect 14875 17728 14887 17731
rect 15930 17728 15936 17740
rect 14875 17700 15936 17728
rect 14875 17697 14887 17700
rect 14829 17691 14887 17697
rect 15930 17688 15936 17700
rect 15988 17688 15994 17740
rect 16209 17731 16267 17737
rect 16209 17697 16221 17731
rect 16255 17728 16267 17731
rect 17681 17731 17739 17737
rect 16255 17700 17632 17728
rect 16255 17697 16267 17700
rect 16209 17691 16267 17697
rect 10994 17632 11652 17660
rect 11698 17620 11704 17672
rect 11756 17660 11762 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 11756 17632 14105 17660
rect 11756 17620 11762 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 15252 17632 15301 17660
rect 15252 17620 15258 17632
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 17604 17660 17632 17700
rect 17681 17697 17693 17731
rect 17727 17728 17739 17731
rect 19904 17728 19932 17768
rect 17727 17700 19932 17728
rect 17727 17697 17739 17700
rect 17681 17691 17739 17697
rect 18693 17663 18751 17669
rect 17604 17632 18644 17660
rect 15289 17623 15347 17629
rect 6822 17592 6828 17604
rect 6564 17564 6828 17592
rect 6822 17552 6828 17564
rect 6880 17552 6886 17604
rect 6932 17564 7314 17592
rect 1765 17527 1823 17533
rect 1765 17493 1777 17527
rect 1811 17524 1823 17527
rect 1946 17524 1952 17536
rect 1811 17496 1952 17524
rect 1811 17493 1823 17496
rect 1765 17487 1823 17493
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 6454 17484 6460 17536
rect 6512 17524 6518 17536
rect 6932 17524 6960 17564
rect 6512 17496 6960 17524
rect 8297 17527 8355 17533
rect 6512 17484 6518 17496
rect 8297 17493 8309 17527
rect 8343 17524 8355 17527
rect 8662 17524 8668 17536
rect 8343 17496 8668 17524
rect 8343 17493 8355 17496
rect 8297 17487 8355 17493
rect 8662 17484 8668 17496
rect 8720 17484 8726 17536
rect 9600 17524 9628 17620
rect 9766 17552 9772 17604
rect 9824 17592 9830 17604
rect 9861 17595 9919 17601
rect 9861 17592 9873 17595
rect 9824 17564 9873 17592
rect 9824 17552 9830 17564
rect 9861 17561 9873 17564
rect 9907 17561 9919 17595
rect 11790 17592 11796 17604
rect 11751 17564 11796 17592
rect 9861 17555 9919 17561
rect 11790 17552 11796 17564
rect 11848 17552 11854 17604
rect 18414 17592 18420 17604
rect 17434 17564 18420 17592
rect 18414 17552 18420 17564
rect 18472 17552 18478 17604
rect 18616 17592 18644 17632
rect 18693 17629 18705 17663
rect 18739 17660 18751 17663
rect 19794 17660 19800 17672
rect 18739 17632 19800 17660
rect 18739 17629 18751 17632
rect 18693 17623 18751 17629
rect 19794 17620 19800 17632
rect 19852 17620 19858 17672
rect 19889 17663 19947 17669
rect 19889 17629 19901 17663
rect 19935 17629 19947 17663
rect 20438 17660 20444 17672
rect 20399 17632 20444 17660
rect 19889 17623 19947 17629
rect 19334 17592 19340 17604
rect 18616 17564 19340 17592
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 19904 17592 19932 17623
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 20622 17620 20628 17672
rect 20680 17660 20686 17672
rect 20809 17663 20867 17669
rect 20809 17660 20821 17663
rect 20680 17632 20821 17660
rect 20680 17620 20686 17632
rect 20809 17629 20821 17632
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 21100 17632 22140 17660
rect 20990 17592 20996 17604
rect 19904 17564 20996 17592
rect 20990 17552 20996 17564
rect 21048 17552 21054 17604
rect 11882 17524 11888 17536
rect 9600 17496 11888 17524
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 13078 17524 13084 17536
rect 13039 17496 13084 17524
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 15473 17527 15531 17533
rect 15473 17493 15485 17527
rect 15519 17524 15531 17527
rect 17586 17524 17592 17536
rect 15519 17496 17592 17524
rect 15519 17493 15531 17496
rect 15473 17487 15531 17493
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 20438 17484 20444 17536
rect 20496 17524 20502 17536
rect 21100 17524 21128 17632
rect 20496 17496 21128 17524
rect 22112 17524 22140 17632
rect 22370 17620 22376 17672
rect 22428 17660 22434 17672
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 22428 17632 22753 17660
rect 22428 17620 22434 17632
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 22848 17660 22876 17768
rect 23477 17765 23489 17799
rect 23523 17796 23535 17799
rect 24670 17796 24676 17808
rect 23523 17768 24676 17796
rect 23523 17765 23535 17768
rect 23477 17759 23535 17765
rect 24670 17756 24676 17768
rect 24728 17756 24734 17808
rect 30558 17756 30564 17808
rect 30616 17796 30622 17808
rect 31570 17796 31576 17808
rect 30616 17768 31576 17796
rect 30616 17756 30622 17768
rect 31570 17756 31576 17768
rect 31628 17796 31634 17808
rect 31628 17768 31754 17796
rect 31628 17756 31634 17768
rect 23400 17700 28212 17728
rect 23400 17669 23428 17700
rect 23385 17663 23443 17669
rect 23385 17660 23397 17663
rect 22848 17632 23397 17660
rect 22741 17623 22799 17629
rect 23385 17629 23397 17632
rect 23431 17629 23443 17663
rect 25958 17660 25964 17672
rect 23385 17623 23443 17629
rect 23768 17632 25964 17660
rect 22281 17595 22339 17601
rect 22281 17561 22293 17595
rect 22327 17592 22339 17595
rect 23768 17592 23796 17632
rect 25958 17620 25964 17632
rect 26016 17620 26022 17672
rect 26142 17620 26148 17672
rect 26200 17660 26206 17672
rect 28184 17669 28212 17700
rect 28718 17688 28724 17740
rect 28776 17728 28782 17740
rect 28905 17731 28963 17737
rect 28905 17728 28917 17731
rect 28776 17700 28917 17728
rect 28776 17688 28782 17700
rect 28905 17697 28917 17700
rect 28951 17697 28963 17731
rect 31726 17728 31754 17768
rect 37182 17756 37188 17808
rect 37240 17796 37246 17808
rect 42886 17796 42892 17808
rect 37240 17768 42892 17796
rect 37240 17756 37246 17768
rect 42886 17756 42892 17768
rect 42944 17756 42950 17808
rect 51046 17796 51074 17836
rect 52178 17824 52184 17836
rect 52236 17824 52242 17876
rect 52457 17867 52515 17873
rect 52457 17833 52469 17867
rect 52503 17864 52515 17867
rect 53190 17864 53196 17876
rect 52503 17836 53196 17864
rect 52503 17833 52515 17836
rect 52457 17827 52515 17833
rect 53190 17824 53196 17836
rect 53248 17824 53254 17876
rect 53926 17864 53932 17876
rect 53887 17836 53932 17864
rect 53926 17824 53932 17836
rect 53984 17824 53990 17876
rect 54113 17867 54171 17873
rect 54113 17833 54125 17867
rect 54159 17833 54171 17867
rect 54113 17827 54171 17833
rect 54128 17796 54156 17827
rect 56410 17824 56416 17876
rect 56468 17864 56474 17876
rect 58161 17867 58219 17873
rect 58161 17864 58173 17867
rect 56468 17836 58173 17864
rect 56468 17824 56474 17836
rect 58161 17833 58173 17836
rect 58207 17833 58219 17867
rect 58161 17827 58219 17833
rect 48608 17768 51074 17796
rect 53024 17768 54156 17796
rect 32030 17728 32036 17740
rect 31726 17700 32036 17728
rect 28905 17691 28963 17697
rect 32030 17688 32036 17700
rect 32088 17728 32094 17740
rect 33321 17731 33379 17737
rect 33321 17728 33333 17731
rect 32088 17700 33333 17728
rect 32088 17688 32094 17700
rect 33321 17697 33333 17700
rect 33367 17728 33379 17731
rect 34790 17728 34796 17740
rect 33367 17700 34796 17728
rect 33367 17697 33379 17700
rect 33321 17691 33379 17697
rect 34790 17688 34796 17700
rect 34848 17688 34854 17740
rect 36262 17688 36268 17740
rect 36320 17728 36326 17740
rect 37645 17731 37703 17737
rect 37645 17728 37657 17731
rect 36320 17700 37657 17728
rect 36320 17688 36326 17700
rect 37645 17697 37657 17700
rect 37691 17728 37703 17731
rect 38930 17728 38936 17740
rect 37691 17700 38936 17728
rect 37691 17697 37703 17700
rect 37645 17691 37703 17697
rect 38930 17688 38936 17700
rect 38988 17688 38994 17740
rect 40405 17731 40463 17737
rect 40405 17697 40417 17731
rect 40451 17728 40463 17731
rect 41598 17728 41604 17740
rect 40451 17700 41604 17728
rect 40451 17697 40463 17700
rect 40405 17691 40463 17697
rect 41598 17688 41604 17700
rect 41656 17688 41662 17740
rect 43806 17728 43812 17740
rect 43767 17700 43812 17728
rect 43806 17688 43812 17700
rect 43864 17688 43870 17740
rect 47394 17728 47400 17740
rect 44192 17700 47400 17728
rect 44192 17672 44220 17700
rect 47394 17688 47400 17700
rect 47452 17688 47458 17740
rect 47581 17731 47639 17737
rect 47581 17697 47593 17731
rect 47627 17728 47639 17731
rect 47670 17728 47676 17740
rect 47627 17700 47676 17728
rect 47627 17697 47639 17700
rect 47581 17691 47639 17697
rect 47670 17688 47676 17700
rect 47728 17688 47734 17740
rect 47857 17731 47915 17737
rect 47857 17697 47869 17731
rect 47903 17728 47915 17731
rect 48038 17728 48044 17740
rect 47903 17700 48044 17728
rect 47903 17697 47915 17700
rect 47857 17691 47915 17697
rect 48038 17688 48044 17700
rect 48096 17688 48102 17740
rect 48608 17737 48636 17768
rect 48593 17731 48651 17737
rect 48593 17728 48605 17731
rect 48240 17700 48605 17728
rect 27985 17663 28043 17669
rect 27985 17660 27997 17663
rect 26200 17632 27997 17660
rect 26200 17620 26206 17632
rect 27985 17629 27997 17632
rect 28031 17629 28043 17663
rect 27985 17623 28043 17629
rect 28169 17663 28227 17669
rect 28169 17629 28181 17663
rect 28215 17629 28227 17663
rect 28169 17623 28227 17629
rect 31662 17620 31668 17672
rect 31720 17660 31726 17672
rect 31757 17663 31815 17669
rect 31757 17660 31769 17663
rect 31720 17632 31769 17660
rect 31720 17620 31726 17632
rect 31757 17629 31769 17632
rect 31803 17629 31815 17663
rect 35250 17660 35256 17672
rect 35211 17632 35256 17660
rect 31757 17623 31815 17629
rect 35250 17620 35256 17632
rect 35308 17620 35314 17672
rect 35894 17660 35900 17672
rect 35855 17632 35900 17660
rect 35894 17620 35900 17632
rect 35952 17620 35958 17672
rect 38102 17660 38108 17672
rect 38063 17632 38108 17660
rect 38102 17620 38108 17632
rect 38160 17620 38166 17672
rect 40310 17660 40316 17672
rect 40271 17632 40316 17660
rect 40310 17620 40316 17632
rect 40368 17620 40374 17672
rect 40957 17663 41015 17669
rect 40957 17629 40969 17663
rect 41003 17660 41015 17663
rect 41003 17632 41184 17660
rect 41003 17629 41015 17632
rect 40957 17623 41015 17629
rect 22327 17564 23796 17592
rect 22327 17561 22339 17564
rect 22281 17555 22339 17561
rect 23842 17552 23848 17604
rect 23900 17592 23906 17604
rect 24949 17595 25007 17601
rect 24949 17592 24961 17595
rect 23900 17564 24961 17592
rect 23900 17552 23906 17564
rect 24949 17561 24961 17564
rect 24995 17561 25007 17595
rect 24949 17555 25007 17561
rect 27338 17552 27344 17604
rect 27396 17592 27402 17604
rect 27433 17595 27491 17601
rect 27433 17592 27445 17595
rect 27396 17564 27445 17592
rect 27396 17552 27402 17564
rect 27433 17561 27445 17564
rect 27479 17592 27491 17595
rect 31202 17592 31208 17604
rect 27479 17564 29868 17592
rect 31163 17564 31208 17592
rect 27479 17561 27491 17564
rect 27433 17555 27491 17561
rect 24397 17527 24455 17533
rect 24397 17524 24409 17527
rect 22112 17496 24409 17524
rect 20496 17484 20502 17496
rect 24397 17493 24409 17496
rect 24443 17493 24455 17527
rect 24397 17487 24455 17493
rect 29641 17527 29699 17533
rect 29641 17493 29653 17527
rect 29687 17524 29699 17527
rect 29730 17524 29736 17536
rect 29687 17496 29736 17524
rect 29687 17493 29699 17496
rect 29641 17487 29699 17493
rect 29730 17484 29736 17496
rect 29788 17484 29794 17536
rect 29840 17524 29868 17564
rect 31202 17552 31208 17564
rect 31260 17592 31266 17604
rect 31941 17595 31999 17601
rect 31941 17592 31953 17595
rect 31260 17564 31953 17592
rect 31260 17552 31266 17564
rect 31941 17561 31953 17564
rect 31987 17561 31999 17595
rect 31941 17555 31999 17561
rect 32306 17552 32312 17604
rect 32364 17592 32370 17604
rect 35802 17592 35808 17604
rect 32364 17564 35808 17592
rect 32364 17552 32370 17564
rect 35802 17552 35808 17564
rect 35860 17552 35866 17604
rect 36170 17592 36176 17604
rect 36131 17564 36176 17592
rect 36170 17552 36176 17564
rect 36228 17552 36234 17604
rect 38838 17592 38844 17604
rect 37398 17564 38844 17592
rect 33318 17524 33324 17536
rect 29840 17496 33324 17524
rect 33318 17484 33324 17496
rect 33376 17484 33382 17536
rect 34054 17524 34060 17536
rect 34015 17496 34060 17524
rect 34054 17484 34060 17496
rect 34112 17524 34118 17536
rect 34606 17524 34612 17536
rect 34112 17496 34612 17524
rect 34112 17484 34118 17496
rect 34606 17484 34612 17496
rect 34664 17484 34670 17536
rect 35345 17527 35403 17533
rect 35345 17493 35357 17527
rect 35391 17524 35403 17527
rect 37476 17524 37504 17564
rect 38838 17552 38844 17564
rect 38896 17552 38902 17604
rect 39114 17592 39120 17604
rect 39075 17564 39120 17592
rect 39114 17552 39120 17564
rect 39172 17552 39178 17604
rect 39301 17595 39359 17601
rect 39301 17561 39313 17595
rect 39347 17592 39359 17595
rect 41156 17592 41184 17632
rect 41230 17620 41236 17672
rect 41288 17660 41294 17672
rect 41417 17663 41475 17669
rect 41417 17660 41429 17663
rect 41288 17632 41429 17660
rect 41288 17620 41294 17632
rect 41417 17629 41429 17632
rect 41463 17660 41475 17663
rect 42058 17660 42064 17672
rect 41463 17632 42064 17660
rect 41463 17629 41475 17632
rect 41417 17623 41475 17629
rect 42058 17620 42064 17632
rect 42116 17620 42122 17672
rect 44174 17660 44180 17672
rect 44135 17632 44180 17660
rect 44174 17620 44180 17632
rect 44232 17620 44238 17672
rect 45002 17660 45008 17672
rect 44963 17632 45008 17660
rect 45002 17620 45008 17632
rect 45060 17620 45066 17672
rect 47489 17663 47547 17669
rect 47489 17629 47501 17663
rect 47535 17660 47547 17663
rect 48240 17660 48268 17700
rect 48593 17697 48605 17700
rect 48639 17697 48651 17731
rect 50430 17728 50436 17740
rect 50391 17700 50436 17728
rect 48593 17691 48651 17697
rect 50430 17688 50436 17700
rect 50488 17688 50494 17740
rect 52362 17728 52368 17740
rect 51046 17700 52368 17728
rect 47535 17632 48268 17660
rect 47535 17629 47547 17632
rect 47489 17623 47547 17629
rect 48314 17620 48320 17672
rect 48372 17660 48378 17672
rect 48372 17632 48417 17660
rect 48372 17620 48378 17632
rect 49050 17620 49056 17672
rect 49108 17660 49114 17672
rect 50341 17663 50399 17669
rect 50341 17660 50353 17663
rect 49108 17632 50353 17660
rect 49108 17620 49114 17632
rect 50341 17629 50353 17632
rect 50387 17660 50399 17663
rect 51046 17660 51074 17700
rect 52362 17688 52368 17700
rect 52420 17728 52426 17740
rect 53024 17728 53052 17768
rect 52420 17700 53052 17728
rect 52420 17688 52426 17700
rect 50387 17632 51074 17660
rect 51629 17663 51687 17669
rect 50387 17629 50399 17632
rect 50341 17623 50399 17629
rect 51629 17629 51641 17663
rect 51675 17629 51687 17663
rect 51810 17660 51816 17672
rect 51771 17632 51816 17660
rect 51629 17623 51687 17629
rect 39347 17564 41092 17592
rect 41156 17564 42748 17592
rect 39347 17561 39359 17564
rect 39301 17555 39359 17561
rect 35391 17496 37504 17524
rect 35391 17493 35403 17496
rect 35345 17487 35403 17493
rect 38286 17484 38292 17536
rect 38344 17524 38350 17536
rect 40954 17524 40960 17536
rect 38344 17496 40960 17524
rect 38344 17484 38350 17496
rect 40954 17484 40960 17496
rect 41012 17484 41018 17536
rect 41064 17524 41092 17564
rect 41782 17524 41788 17536
rect 41064 17496 41788 17524
rect 41782 17484 41788 17496
rect 41840 17484 41846 17536
rect 42720 17524 42748 17564
rect 42794 17552 42800 17604
rect 42852 17552 42858 17604
rect 45186 17592 45192 17604
rect 45147 17564 45192 17592
rect 45186 17552 45192 17564
rect 45244 17552 45250 17604
rect 45922 17552 45928 17604
rect 45980 17592 45986 17604
rect 46845 17595 46903 17601
rect 46845 17592 46857 17595
rect 45980 17564 46857 17592
rect 45980 17552 45986 17564
rect 46845 17561 46857 17564
rect 46891 17561 46903 17595
rect 46845 17555 46903 17561
rect 49510 17524 49516 17536
rect 42720 17496 49516 17524
rect 49510 17484 49516 17496
rect 49568 17484 49574 17536
rect 51644 17524 51672 17623
rect 51810 17620 51816 17632
rect 51868 17620 51874 17672
rect 52273 17663 52331 17669
rect 52273 17629 52285 17663
rect 52319 17629 52331 17663
rect 52454 17660 52460 17672
rect 52415 17632 52460 17660
rect 52273 17623 52331 17629
rect 51721 17595 51779 17601
rect 51721 17561 51733 17595
rect 51767 17592 51779 17595
rect 52178 17592 52184 17604
rect 51767 17564 52184 17592
rect 51767 17561 51779 17564
rect 51721 17555 51779 17561
rect 52178 17552 52184 17564
rect 52236 17552 52242 17604
rect 52288 17592 52316 17623
rect 52454 17620 52460 17632
rect 52512 17620 52518 17672
rect 52914 17660 52920 17672
rect 52875 17632 52920 17660
rect 52914 17620 52920 17632
rect 52972 17620 52978 17672
rect 53024 17660 53052 17700
rect 54294 17688 54300 17740
rect 54352 17728 54358 17740
rect 55493 17731 55551 17737
rect 55493 17728 55505 17731
rect 54352 17700 55505 17728
rect 54352 17688 54358 17700
rect 55493 17697 55505 17700
rect 55539 17697 55551 17731
rect 55493 17691 55551 17697
rect 56318 17688 56324 17740
rect 56376 17728 56382 17740
rect 56413 17731 56471 17737
rect 56413 17728 56425 17731
rect 56376 17700 56425 17728
rect 56376 17688 56382 17700
rect 56413 17697 56425 17700
rect 56459 17697 56471 17731
rect 56686 17728 56692 17740
rect 56647 17700 56692 17728
rect 56413 17691 56471 17697
rect 56686 17688 56692 17700
rect 56744 17688 56750 17740
rect 54110 17660 54116 17672
rect 53024 17632 53236 17660
rect 54023 17632 54116 17660
rect 52730 17592 52736 17604
rect 52288 17564 52736 17592
rect 52730 17552 52736 17564
rect 52788 17552 52794 17604
rect 53006 17524 53012 17536
rect 51644 17496 53012 17524
rect 53006 17484 53012 17496
rect 53064 17524 53070 17536
rect 53208 17533 53236 17632
rect 54110 17620 54116 17632
rect 54168 17620 54174 17672
rect 54205 17663 54263 17669
rect 54205 17629 54217 17663
rect 54251 17660 54263 17663
rect 54754 17660 54760 17672
rect 54251 17632 54760 17660
rect 54251 17629 54263 17632
rect 54205 17623 54263 17629
rect 54754 17620 54760 17632
rect 54812 17620 54818 17672
rect 55585 17663 55643 17669
rect 55585 17629 55597 17663
rect 55631 17629 55643 17663
rect 55585 17623 55643 17629
rect 53466 17552 53472 17604
rect 53524 17592 53530 17604
rect 53524 17564 53569 17592
rect 53524 17552 53530 17564
rect 53101 17527 53159 17533
rect 53101 17524 53113 17527
rect 53064 17496 53113 17524
rect 53064 17484 53070 17496
rect 53101 17493 53113 17496
rect 53147 17493 53159 17527
rect 53101 17487 53159 17493
rect 53193 17527 53251 17533
rect 53193 17493 53205 17527
rect 53239 17493 53251 17527
rect 53193 17487 53251 17493
rect 53282 17484 53288 17536
rect 53340 17524 53346 17536
rect 54128 17524 54156 17620
rect 54386 17592 54392 17604
rect 54347 17564 54392 17592
rect 54386 17552 54392 17564
rect 54444 17552 54450 17604
rect 55600 17592 55628 17623
rect 56778 17592 56784 17604
rect 55600 17564 56784 17592
rect 55600 17524 55628 17564
rect 56778 17552 56784 17564
rect 56836 17552 56842 17604
rect 57330 17552 57336 17604
rect 57388 17552 57394 17604
rect 53340 17496 53385 17524
rect 54128 17496 55628 17524
rect 55953 17527 56011 17533
rect 53340 17484 53346 17496
rect 55953 17493 55965 17527
rect 55999 17524 56011 17527
rect 56686 17524 56692 17536
rect 55999 17496 56692 17524
rect 55999 17493 56011 17496
rect 55953 17487 56011 17493
rect 56686 17484 56692 17496
rect 56744 17484 56750 17536
rect 1104 17434 58880 17456
rect 1104 17382 15398 17434
rect 15450 17382 15462 17434
rect 15514 17382 15526 17434
rect 15578 17382 15590 17434
rect 15642 17382 15654 17434
rect 15706 17382 29846 17434
rect 29898 17382 29910 17434
rect 29962 17382 29974 17434
rect 30026 17382 30038 17434
rect 30090 17382 30102 17434
rect 30154 17382 44294 17434
rect 44346 17382 44358 17434
rect 44410 17382 44422 17434
rect 44474 17382 44486 17434
rect 44538 17382 44550 17434
rect 44602 17382 58880 17434
rect 1104 17360 58880 17382
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17320 4583 17323
rect 5350 17320 5356 17332
rect 4571 17292 5356 17320
rect 4571 17289 4583 17292
rect 4525 17283 4583 17289
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 5629 17323 5687 17329
rect 5629 17289 5641 17323
rect 5675 17320 5687 17323
rect 7006 17320 7012 17332
rect 5675 17292 7012 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 9125 17323 9183 17329
rect 9125 17320 9137 17323
rect 8628 17292 9137 17320
rect 8628 17280 8634 17292
rect 9125 17289 9137 17292
rect 9171 17289 9183 17323
rect 9125 17283 9183 17289
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 17644 17292 19012 17320
rect 17644 17280 17650 17292
rect 1946 17252 1952 17264
rect 1907 17224 1952 17252
rect 1946 17212 1952 17224
rect 2004 17212 2010 17264
rect 3510 17252 3516 17264
rect 3174 17224 3516 17252
rect 3510 17212 3516 17224
rect 3568 17212 3574 17264
rect 4798 17252 4804 17264
rect 4632 17224 4804 17252
rect 4632 17193 4660 17224
rect 4798 17212 4804 17224
rect 4856 17252 4862 17264
rect 11517 17255 11575 17261
rect 11517 17252 11529 17255
rect 4856 17224 11529 17252
rect 4856 17212 4862 17224
rect 11517 17221 11529 17224
rect 11563 17221 11575 17255
rect 11517 17215 11575 17221
rect 11606 17212 11612 17264
rect 11664 17252 11670 17264
rect 14369 17255 14427 17261
rect 11664 17224 12098 17252
rect 11664 17212 11670 17224
rect 14369 17221 14381 17255
rect 14415 17252 14427 17255
rect 15286 17252 15292 17264
rect 14415 17224 15292 17252
rect 14415 17221 14427 17224
rect 14369 17215 14427 17221
rect 15286 17212 15292 17224
rect 15344 17212 15350 17264
rect 17954 17212 17960 17264
rect 18012 17212 18018 17264
rect 18984 17261 19012 17292
rect 19794 17280 19800 17332
rect 19852 17320 19858 17332
rect 25038 17320 25044 17332
rect 19852 17292 25044 17320
rect 19852 17280 19858 17292
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 25682 17320 25688 17332
rect 25643 17292 25688 17320
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 33965 17323 34023 17329
rect 33965 17320 33977 17323
rect 31496 17292 33977 17320
rect 18969 17255 19027 17261
rect 18969 17221 18981 17255
rect 19015 17221 19027 17255
rect 18969 17215 19027 17221
rect 22922 17212 22928 17264
rect 22980 17252 22986 17264
rect 23569 17255 23627 17261
rect 23569 17252 23581 17255
rect 22980 17224 23581 17252
rect 22980 17212 22986 17224
rect 23569 17221 23581 17224
rect 23615 17221 23627 17255
rect 26329 17255 26387 17261
rect 26329 17252 26341 17255
rect 24794 17224 26341 17252
rect 23569 17215 23627 17221
rect 26329 17221 26341 17224
rect 26375 17221 26387 17255
rect 26329 17215 26387 17221
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17085 1731 17119
rect 1673 17079 1731 17085
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17085 3755 17119
rect 3697 17079 3755 17085
rect 1688 16980 1716 17079
rect 3050 17008 3056 17060
rect 3108 17048 3114 17060
rect 3712 17048 3740 17079
rect 5276 17060 5304 17147
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 6546 17184 6552 17196
rect 5960 17156 6552 17184
rect 5960 17144 5966 17156
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17184 7895 17187
rect 9122 17184 9128 17196
rect 7883 17156 9128 17184
rect 7883 17153 7895 17156
rect 7837 17147 7895 17153
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 10318 17184 10324 17196
rect 10279 17156 10324 17184
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 10778 17184 10784 17196
rect 10739 17156 10784 17184
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 16540 17156 16681 17184
rect 16540 17144 16546 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 18432 17156 21772 17184
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17116 5411 17119
rect 5442 17116 5448 17128
rect 5399 17088 5448 17116
rect 5399 17085 5411 17088
rect 5353 17079 5411 17085
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 6730 17116 6736 17128
rect 6687 17088 6736 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 6730 17076 6736 17088
rect 6788 17076 6794 17128
rect 8754 17116 8760 17128
rect 6840 17088 8760 17116
rect 5258 17048 5264 17060
rect 3108 17020 3740 17048
rect 5171 17020 5264 17048
rect 3108 17008 3114 17020
rect 5258 17008 5264 17020
rect 5316 17048 5322 17060
rect 6840 17048 6868 17088
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 11112 17088 13277 17116
rect 11112 17076 11118 17088
rect 13265 17085 13277 17088
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 16574 17116 16580 17128
rect 13587 17088 16580 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 17954 17116 17960 17128
rect 16991 17088 17960 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 18432 17125 18460 17156
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17085 18475 17119
rect 20714 17116 20720 17128
rect 20675 17088 20720 17116
rect 18417 17079 18475 17085
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 5316 17020 6868 17048
rect 6917 17051 6975 17057
rect 5316 17008 5322 17020
rect 6917 17017 6929 17051
rect 6963 17048 6975 17051
rect 7374 17048 7380 17060
rect 6963 17020 7380 17048
rect 6963 17017 6975 17020
rect 6917 17011 6975 17017
rect 7374 17008 7380 17020
rect 7432 17008 7438 17060
rect 10229 17051 10287 17057
rect 10229 17017 10241 17051
rect 10275 17048 10287 17051
rect 12250 17048 12256 17060
rect 10275 17020 12256 17048
rect 10275 17017 10287 17020
rect 10229 17011 10287 17017
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 21174 17048 21180 17060
rect 21135 17020 21180 17048
rect 21174 17008 21180 17020
rect 21232 17008 21238 17060
rect 21744 17048 21772 17156
rect 21818 17144 21824 17196
rect 21876 17182 21882 17196
rect 22657 17185 22715 17191
rect 21876 17154 21919 17182
rect 21876 17144 21882 17154
rect 22657 17151 22669 17185
rect 22703 17182 22715 17185
rect 23290 17184 23296 17196
rect 22703 17174 22784 17182
rect 22703 17154 22876 17174
rect 23251 17156 23296 17184
rect 22703 17151 22715 17154
rect 22657 17145 22715 17151
rect 22756 17146 22876 17154
rect 22848 17116 22876 17146
rect 23290 17144 23296 17156
rect 23348 17144 23354 17196
rect 24854 17144 24860 17196
rect 24912 17184 24918 17196
rect 25777 17187 25835 17193
rect 25777 17184 25789 17187
rect 24912 17156 25789 17184
rect 24912 17144 24918 17156
rect 25777 17153 25789 17156
rect 25823 17184 25835 17187
rect 26237 17187 26295 17193
rect 26237 17184 26249 17187
rect 25823 17156 26249 17184
rect 25823 17153 25835 17156
rect 25777 17147 25835 17153
rect 26237 17153 26249 17156
rect 26283 17153 26295 17187
rect 26237 17147 26295 17153
rect 28074 17144 28080 17196
rect 28132 17184 28138 17196
rect 28169 17187 28227 17193
rect 28169 17184 28181 17187
rect 28132 17156 28181 17184
rect 28132 17144 28138 17156
rect 28169 17153 28181 17156
rect 28215 17153 28227 17187
rect 28350 17184 28356 17196
rect 28311 17156 28356 17184
rect 28169 17147 28227 17153
rect 28350 17144 28356 17156
rect 28408 17144 28414 17196
rect 30009 17187 30067 17193
rect 30009 17153 30021 17187
rect 30055 17184 30067 17187
rect 31386 17184 31392 17196
rect 30055 17156 31392 17184
rect 30055 17153 30067 17156
rect 30009 17147 30067 17153
rect 31386 17144 31392 17156
rect 31444 17144 31450 17196
rect 31496 17193 31524 17292
rect 33965 17289 33977 17292
rect 34011 17320 34023 17323
rect 35529 17323 35587 17329
rect 34011 17292 35020 17320
rect 34011 17289 34023 17292
rect 33965 17283 34023 17289
rect 32582 17252 32588 17264
rect 31588 17224 32588 17252
rect 31481 17187 31539 17193
rect 31481 17153 31493 17187
rect 31527 17153 31539 17187
rect 31481 17147 31539 17153
rect 24946 17116 24952 17128
rect 22848 17088 24952 17116
rect 22848 17048 22876 17088
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 29178 17116 29184 17128
rect 29139 17088 29184 17116
rect 29178 17076 29184 17088
rect 29236 17076 29242 17128
rect 29270 17076 29276 17128
rect 29328 17116 29334 17128
rect 29917 17119 29975 17125
rect 29917 17116 29929 17119
rect 29328 17088 29929 17116
rect 29328 17076 29334 17088
rect 29917 17085 29929 17088
rect 29963 17085 29975 17119
rect 29917 17079 29975 17085
rect 30098 17076 30104 17128
rect 30156 17116 30162 17128
rect 31588 17116 31616 17224
rect 32582 17212 32588 17224
rect 32640 17212 32646 17264
rect 34790 17252 34796 17264
rect 33718 17224 34796 17252
rect 34790 17212 34796 17224
rect 34848 17212 34854 17264
rect 34698 17184 34704 17196
rect 34659 17156 34704 17184
rect 34698 17144 34704 17156
rect 34756 17144 34762 17196
rect 34992 17193 35020 17292
rect 35529 17289 35541 17323
rect 35575 17320 35587 17323
rect 37182 17320 37188 17332
rect 35575 17292 37188 17320
rect 35575 17289 35587 17292
rect 35529 17283 35587 17289
rect 37182 17280 37188 17292
rect 37240 17280 37246 17332
rect 38562 17320 38568 17332
rect 37936 17292 38568 17320
rect 35802 17212 35808 17264
rect 35860 17252 35866 17264
rect 37936 17252 37964 17292
rect 38562 17280 38568 17292
rect 38620 17280 38626 17332
rect 41877 17323 41935 17329
rect 41877 17289 41889 17323
rect 41923 17320 41935 17323
rect 44174 17320 44180 17332
rect 41923 17292 44180 17320
rect 41923 17289 41935 17292
rect 41877 17283 41935 17289
rect 44174 17280 44180 17292
rect 44232 17280 44238 17332
rect 44818 17280 44824 17332
rect 44876 17320 44882 17332
rect 44876 17292 45416 17320
rect 44876 17280 44882 17292
rect 38838 17252 38844 17264
rect 35860 17224 37964 17252
rect 38778 17224 38844 17252
rect 35860 17212 35866 17224
rect 38838 17212 38844 17224
rect 38896 17212 38902 17264
rect 40770 17212 40776 17264
rect 40828 17212 40834 17264
rect 45388 17261 45416 17292
rect 46750 17280 46756 17332
rect 46808 17320 46814 17332
rect 47581 17323 47639 17329
rect 47581 17320 47593 17323
rect 46808 17292 47593 17320
rect 46808 17280 46814 17292
rect 47581 17289 47593 17292
rect 47627 17289 47639 17323
rect 48590 17320 48596 17332
rect 48551 17292 48596 17320
rect 47581 17283 47639 17289
rect 48590 17280 48596 17292
rect 48648 17280 48654 17332
rect 51810 17280 51816 17332
rect 51868 17320 51874 17332
rect 53466 17320 53472 17332
rect 51868 17292 53472 17320
rect 51868 17280 51874 17292
rect 53466 17280 53472 17292
rect 53524 17280 53530 17332
rect 53558 17280 53564 17332
rect 53616 17320 53622 17332
rect 55125 17323 55183 17329
rect 55125 17320 55137 17323
rect 53616 17292 55137 17320
rect 53616 17280 53622 17292
rect 55125 17289 55137 17292
rect 55171 17289 55183 17323
rect 55125 17283 55183 17289
rect 55493 17323 55551 17329
rect 55493 17289 55505 17323
rect 55539 17320 55551 17323
rect 56226 17320 56232 17332
rect 55539 17292 56232 17320
rect 55539 17289 55551 17292
rect 55493 17283 55551 17289
rect 56226 17280 56232 17292
rect 56284 17280 56290 17332
rect 57882 17320 57888 17332
rect 57843 17292 57888 17320
rect 57882 17280 57888 17292
rect 57940 17280 57946 17332
rect 45373 17255 45431 17261
rect 45373 17221 45385 17255
rect 45419 17221 45431 17255
rect 49050 17252 49056 17264
rect 45373 17215 45431 17221
rect 47596 17224 49056 17252
rect 34977 17187 35035 17193
rect 34977 17153 34989 17187
rect 35023 17153 35035 17187
rect 34977 17147 35035 17153
rect 36265 17187 36323 17193
rect 36265 17153 36277 17187
rect 36311 17184 36323 17187
rect 36446 17184 36452 17196
rect 36311 17156 36452 17184
rect 36311 17153 36323 17156
rect 36265 17147 36323 17153
rect 36446 17144 36452 17156
rect 36504 17144 36510 17196
rect 39482 17184 39488 17196
rect 39443 17156 39488 17184
rect 39482 17144 39488 17156
rect 39540 17144 39546 17196
rect 41693 17187 41751 17193
rect 41693 17153 41705 17187
rect 41739 17184 41751 17187
rect 41782 17184 41788 17196
rect 41739 17156 41788 17184
rect 41739 17153 41751 17156
rect 41693 17147 41751 17153
rect 41782 17144 41788 17156
rect 41840 17144 41846 17196
rect 32214 17116 32220 17128
rect 30156 17088 31616 17116
rect 32175 17088 32220 17116
rect 30156 17076 30162 17088
rect 32214 17076 32220 17088
rect 32272 17076 32278 17128
rect 32493 17119 32551 17125
rect 32493 17085 32505 17119
rect 32539 17116 32551 17119
rect 33226 17116 33232 17128
rect 32539 17088 33232 17116
rect 32539 17085 32551 17088
rect 32493 17079 32551 17085
rect 33226 17076 33232 17088
rect 33284 17076 33290 17128
rect 35986 17076 35992 17128
rect 36044 17116 36050 17128
rect 37277 17119 37335 17125
rect 37277 17116 37289 17119
rect 36044 17088 37289 17116
rect 36044 17076 36050 17088
rect 37277 17085 37289 17088
rect 37323 17085 37335 17119
rect 37277 17079 37335 17085
rect 37553 17119 37611 17125
rect 37553 17085 37565 17119
rect 37599 17116 37611 17119
rect 38562 17116 38568 17128
rect 37599 17088 38568 17116
rect 37599 17085 37611 17088
rect 37553 17079 37611 17085
rect 38562 17076 38568 17088
rect 38620 17076 38626 17128
rect 39758 17116 39764 17128
rect 39719 17088 39764 17116
rect 39758 17076 39764 17088
rect 39816 17076 39822 17128
rect 42613 17119 42671 17125
rect 42613 17085 42625 17119
rect 42659 17085 42671 17119
rect 42613 17079 42671 17085
rect 21744 17020 22876 17048
rect 27617 17051 27675 17057
rect 27617 17017 27629 17051
rect 27663 17048 27675 17051
rect 28810 17048 28816 17060
rect 27663 17020 28816 17048
rect 27663 17017 27675 17020
rect 27617 17011 27675 17017
rect 28810 17008 28816 17020
rect 28868 17008 28874 17060
rect 29638 17048 29644 17060
rect 29599 17020 29644 17048
rect 29638 17008 29644 17020
rect 29696 17008 29702 17060
rect 36354 17048 36360 17060
rect 33520 17020 36360 17048
rect 3142 16980 3148 16992
rect 1688 16952 3148 16980
rect 3142 16940 3148 16952
rect 3200 16980 3206 16992
rect 3418 16980 3424 16992
rect 3200 16952 3424 16980
rect 3200 16940 3206 16952
rect 3418 16940 3424 16952
rect 3476 16940 3482 16992
rect 10873 16983 10931 16989
rect 10873 16949 10885 16983
rect 10919 16980 10931 16983
rect 12710 16980 12716 16992
rect 10919 16952 12716 16980
rect 10919 16949 10931 16952
rect 10873 16943 10931 16949
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 15841 16983 15899 16989
rect 15841 16949 15853 16983
rect 15887 16980 15899 16983
rect 18230 16980 18236 16992
rect 15887 16952 18236 16980
rect 15887 16949 15899 16952
rect 15841 16943 15899 16949
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 21913 16983 21971 16989
rect 21913 16949 21925 16983
rect 21959 16980 21971 16983
rect 22278 16980 22284 16992
rect 21959 16952 22284 16980
rect 21959 16949 21971 16952
rect 21913 16943 21971 16949
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 22741 16983 22799 16989
rect 22741 16949 22753 16983
rect 22787 16980 22799 16983
rect 23198 16980 23204 16992
rect 22787 16952 23204 16980
rect 22787 16949 22799 16952
rect 22741 16943 22799 16949
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 25038 16940 25044 16992
rect 25096 16980 25102 16992
rect 26418 16980 26424 16992
rect 25096 16952 26424 16980
rect 25096 16940 25102 16952
rect 26418 16940 26424 16952
rect 26476 16940 26482 16992
rect 26970 16980 26976 16992
rect 26931 16952 26976 16980
rect 26970 16940 26976 16952
rect 27028 16940 27034 16992
rect 30745 16983 30803 16989
rect 30745 16949 30757 16983
rect 30791 16980 30803 16983
rect 31018 16980 31024 16992
rect 30791 16952 31024 16980
rect 30791 16949 30803 16952
rect 30745 16943 30803 16949
rect 31018 16940 31024 16952
rect 31076 16940 31082 16992
rect 31294 16980 31300 16992
rect 31255 16952 31300 16980
rect 31294 16940 31300 16952
rect 31352 16940 31358 16992
rect 32582 16940 32588 16992
rect 32640 16980 32646 16992
rect 33520 16980 33548 17020
rect 36354 17008 36360 17020
rect 36412 17008 36418 17060
rect 42628 17048 42656 17079
rect 42886 17076 42892 17128
rect 42944 17116 42950 17128
rect 44085 17119 44143 17125
rect 44085 17116 44097 17119
rect 42944 17088 44097 17116
rect 42944 17076 42950 17088
rect 44085 17085 44097 17088
rect 44131 17085 44143 17119
rect 44085 17079 44143 17085
rect 44269 17119 44327 17125
rect 44269 17085 44281 17119
rect 44315 17085 44327 17119
rect 44269 17079 44327 17085
rect 45189 17119 45247 17125
rect 45189 17085 45201 17119
rect 45235 17116 45247 17119
rect 45646 17116 45652 17128
rect 45235 17088 45652 17116
rect 45235 17085 45247 17088
rect 45189 17079 45247 17085
rect 43530 17048 43536 17060
rect 42628 17020 43536 17048
rect 43530 17008 43536 17020
rect 43588 17008 43594 17060
rect 44284 17048 44312 17079
rect 45646 17076 45652 17088
rect 45704 17076 45710 17128
rect 45922 17116 45928 17128
rect 45883 17088 45928 17116
rect 45922 17076 45928 17088
rect 45980 17076 45986 17128
rect 47596 17048 47624 17224
rect 49050 17212 49056 17224
rect 49108 17212 49114 17264
rect 49786 17252 49792 17264
rect 49436 17224 49792 17252
rect 47762 17184 47768 17196
rect 47723 17156 47768 17184
rect 47762 17144 47768 17156
rect 47820 17144 47826 17196
rect 47857 17187 47915 17193
rect 47857 17153 47869 17187
rect 47903 17153 47915 17187
rect 48038 17184 48044 17196
rect 47999 17156 48044 17184
rect 47857 17147 47915 17153
rect 47872 17116 47900 17147
rect 48038 17144 48044 17156
rect 48096 17144 48102 17196
rect 49436 17193 49464 17224
rect 49786 17212 49792 17224
rect 49844 17212 49850 17264
rect 50246 17212 50252 17264
rect 50304 17212 50310 17264
rect 52914 17212 52920 17264
rect 52972 17252 52978 17264
rect 55950 17252 55956 17264
rect 52972 17224 53017 17252
rect 55911 17224 55956 17252
rect 52972 17212 52978 17224
rect 55950 17212 55956 17224
rect 56008 17212 56014 17264
rect 48133 17187 48191 17193
rect 48133 17153 48145 17187
rect 48179 17184 48191 17187
rect 49421 17187 49479 17193
rect 48179 17156 48268 17184
rect 48179 17153 48191 17156
rect 48133 17147 48191 17153
rect 47872 17088 48176 17116
rect 48148 17060 48176 17088
rect 44284 17020 47624 17048
rect 48130 17008 48136 17060
rect 48188 17008 48194 17060
rect 36078 16980 36084 16992
rect 32640 16952 33548 16980
rect 36039 16952 36084 16980
rect 32640 16940 32646 16952
rect 36078 16940 36084 16952
rect 36136 16980 36142 16992
rect 38286 16980 38292 16992
rect 36136 16952 38292 16980
rect 36136 16940 36142 16952
rect 38286 16940 38292 16952
rect 38344 16940 38350 16992
rect 39022 16980 39028 16992
rect 38983 16952 39028 16980
rect 39022 16940 39028 16952
rect 39080 16940 39086 16992
rect 41230 16980 41236 16992
rect 41191 16952 41236 16980
rect 41230 16940 41236 16952
rect 41288 16940 41294 16992
rect 47670 16940 47676 16992
rect 47728 16980 47734 16992
rect 48240 16980 48268 17156
rect 49421 17153 49433 17187
rect 49467 17153 49479 17187
rect 51902 17184 51908 17196
rect 51863 17156 51908 17184
rect 49421 17147 49479 17153
rect 51902 17144 51908 17156
rect 51960 17144 51966 17196
rect 52181 17187 52239 17193
rect 52181 17153 52193 17187
rect 52227 17184 52239 17187
rect 52546 17184 52552 17196
rect 52227 17156 52552 17184
rect 52227 17153 52239 17156
rect 52181 17147 52239 17153
rect 52546 17144 52552 17156
rect 52604 17144 52610 17196
rect 52730 17184 52736 17196
rect 52691 17156 52736 17184
rect 52730 17144 52736 17156
rect 52788 17144 52794 17196
rect 55030 17184 55036 17196
rect 54991 17156 55036 17184
rect 55030 17144 55036 17156
rect 55088 17144 55094 17196
rect 55214 17144 55220 17196
rect 55272 17184 55278 17196
rect 55309 17187 55367 17193
rect 55309 17184 55321 17187
rect 55272 17156 55321 17184
rect 55272 17144 55278 17156
rect 55309 17153 55321 17156
rect 55355 17153 55367 17187
rect 58069 17187 58127 17193
rect 58069 17184 58081 17187
rect 55309 17147 55367 17153
rect 57256 17156 58081 17184
rect 49697 17119 49755 17125
rect 49697 17085 49709 17119
rect 49743 17116 49755 17119
rect 50154 17116 50160 17128
rect 49743 17088 50160 17116
rect 49743 17085 49755 17088
rect 49697 17079 49755 17085
rect 50154 17076 50160 17088
rect 50212 17076 50218 17128
rect 52089 17119 52147 17125
rect 52089 17085 52101 17119
rect 52135 17116 52147 17119
rect 52362 17116 52368 17128
rect 52135 17088 52368 17116
rect 52135 17085 52147 17088
rect 52089 17079 52147 17085
rect 52362 17076 52368 17088
rect 52420 17076 52426 17128
rect 54202 17116 54208 17128
rect 54163 17088 54208 17116
rect 54202 17076 54208 17088
rect 54260 17076 54266 17128
rect 57256 17060 57284 17156
rect 58069 17153 58081 17156
rect 58115 17153 58127 17187
rect 58069 17147 58127 17153
rect 51169 17051 51227 17057
rect 51169 17017 51181 17051
rect 51215 17048 51227 17051
rect 51442 17048 51448 17060
rect 51215 17020 51448 17048
rect 51215 17017 51227 17020
rect 51169 17011 51227 17017
rect 51442 17008 51448 17020
rect 51500 17048 51506 17060
rect 51500 17020 51948 17048
rect 51500 17008 51506 17020
rect 47728 16952 48268 16980
rect 47728 16940 47734 16952
rect 51350 16940 51356 16992
rect 51408 16980 51414 16992
rect 51920 16989 51948 17020
rect 52178 17008 52184 17060
rect 52236 17048 52242 17060
rect 53926 17048 53932 17060
rect 52236 17020 53932 17048
rect 52236 17008 52242 17020
rect 53926 17008 53932 17020
rect 53984 17008 53990 17060
rect 57238 17048 57244 17060
rect 57199 17020 57244 17048
rect 57238 17008 57244 17020
rect 57296 17008 57302 17060
rect 51721 16983 51779 16989
rect 51721 16980 51733 16983
rect 51408 16952 51733 16980
rect 51408 16940 51414 16952
rect 51721 16949 51733 16952
rect 51767 16949 51779 16983
rect 51721 16943 51779 16949
rect 51905 16983 51963 16989
rect 51905 16949 51917 16983
rect 51951 16949 51963 16983
rect 51905 16943 51963 16949
rect 52546 16940 52552 16992
rect 52604 16980 52610 16992
rect 52730 16980 52736 16992
rect 52604 16952 52736 16980
rect 52604 16940 52610 16952
rect 52730 16940 52736 16952
rect 52788 16980 52794 16992
rect 53190 16980 53196 16992
rect 52788 16952 53196 16980
rect 52788 16940 52794 16952
rect 53190 16940 53196 16952
rect 53248 16940 53254 16992
rect 1104 16890 58880 16912
rect 1104 16838 8174 16890
rect 8226 16838 8238 16890
rect 8290 16838 8302 16890
rect 8354 16838 8366 16890
rect 8418 16838 8430 16890
rect 8482 16838 22622 16890
rect 22674 16838 22686 16890
rect 22738 16838 22750 16890
rect 22802 16838 22814 16890
rect 22866 16838 22878 16890
rect 22930 16838 37070 16890
rect 37122 16838 37134 16890
rect 37186 16838 37198 16890
rect 37250 16838 37262 16890
rect 37314 16838 37326 16890
rect 37378 16838 51518 16890
rect 51570 16838 51582 16890
rect 51634 16838 51646 16890
rect 51698 16838 51710 16890
rect 51762 16838 51774 16890
rect 51826 16838 58880 16890
rect 1104 16816 58880 16838
rect 6086 16776 6092 16788
rect 3988 16748 6092 16776
rect 3237 16643 3295 16649
rect 3237 16609 3249 16643
rect 3283 16640 3295 16643
rect 3283 16612 3740 16640
rect 3283 16609 3295 16612
rect 3237 16603 3295 16609
rect 3712 16504 3740 16612
rect 3878 16572 3884 16584
rect 3839 16544 3884 16572
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 3988 16581 4016 16748
rect 6086 16736 6092 16748
rect 6144 16736 6150 16788
rect 8036 16748 9168 16776
rect 8036 16708 8064 16748
rect 9030 16708 9036 16720
rect 4632 16680 8064 16708
rect 8404 16680 9036 16708
rect 4632 16581 4660 16680
rect 6270 16640 6276 16652
rect 6231 16612 6276 16640
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 8404 16649 8432 16680
rect 9030 16668 9036 16680
rect 9088 16668 9094 16720
rect 9140 16708 9168 16748
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 17770 16776 17776 16788
rect 16632 16748 17776 16776
rect 16632 16736 16638 16748
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 17862 16736 17868 16788
rect 17920 16776 17926 16788
rect 21637 16779 21695 16785
rect 17920 16748 21588 16776
rect 17920 16736 17926 16748
rect 13262 16708 13268 16720
rect 9140 16680 9536 16708
rect 13175 16680 13268 16708
rect 9508 16652 9536 16680
rect 6733 16643 6791 16649
rect 6733 16640 6745 16643
rect 6604 16612 6745 16640
rect 6604 16600 6610 16612
rect 6733 16609 6745 16612
rect 6779 16609 6791 16643
rect 6733 16603 6791 16609
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8389 16643 8447 16649
rect 7883 16612 8340 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 5166 16572 5172 16584
rect 5127 16544 5172 16572
rect 4617 16535 4675 16541
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5261 16575 5319 16581
rect 5261 16541 5273 16575
rect 5307 16572 5319 16575
rect 5442 16572 5448 16584
rect 5307 16544 5448 16572
rect 5307 16541 5319 16544
rect 5261 16535 5319 16541
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 6181 16575 6239 16581
rect 6181 16541 6193 16575
rect 6227 16572 6239 16575
rect 7190 16572 7196 16584
rect 6227 16544 7196 16572
rect 6227 16541 6239 16544
rect 6181 16535 6239 16541
rect 7190 16532 7196 16544
rect 7248 16532 7254 16584
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16541 7619 16575
rect 8312 16572 8340 16612
rect 8389 16609 8401 16643
rect 8435 16609 8447 16643
rect 9490 16640 9496 16652
rect 9451 16612 9496 16640
rect 8389 16603 8447 16609
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 10778 16600 10784 16652
rect 10836 16640 10842 16652
rect 10836 16612 10916 16640
rect 10836 16600 10842 16612
rect 8754 16572 8760 16584
rect 8312 16544 8760 16572
rect 7561 16535 7619 16541
rect 5350 16504 5356 16516
rect 3712 16476 5356 16504
rect 5350 16464 5356 16476
rect 5408 16464 5414 16516
rect 5534 16464 5540 16516
rect 5592 16504 5598 16516
rect 6362 16504 6368 16516
rect 5592 16476 6368 16504
rect 5592 16464 5598 16476
rect 6362 16464 6368 16476
rect 6420 16504 6426 16516
rect 7576 16504 7604 16535
rect 8754 16532 8760 16544
rect 8812 16532 8818 16584
rect 9214 16572 9220 16584
rect 9175 16544 9220 16572
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 10888 16581 10916 16612
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 13188 16649 13216 16680
rect 13262 16668 13268 16680
rect 13320 16708 13326 16720
rect 16482 16708 16488 16720
rect 13320 16680 16488 16708
rect 13320 16668 13326 16680
rect 16482 16668 16488 16680
rect 16540 16668 16546 16720
rect 19334 16708 19340 16720
rect 18156 16680 19340 16708
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 11296 16612 12909 16640
rect 11296 16600 11302 16612
rect 12897 16609 12909 16612
rect 12943 16609 12955 16643
rect 12897 16603 12955 16609
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 14826 16600 14832 16652
rect 14884 16640 14890 16652
rect 15010 16640 15016 16652
rect 14884 16612 15016 16640
rect 14884 16600 14890 16612
rect 14936 16581 14964 16612
rect 15010 16600 15016 16612
rect 15068 16600 15074 16652
rect 16574 16640 16580 16652
rect 15396 16612 16580 16640
rect 15396 16581 15424 16612
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16640 17647 16643
rect 18156 16640 18184 16680
rect 19334 16668 19340 16680
rect 19392 16668 19398 16720
rect 21560 16708 21588 16748
rect 21637 16745 21649 16779
rect 21683 16776 21695 16779
rect 23014 16776 23020 16788
rect 21683 16748 23020 16776
rect 21683 16745 21695 16748
rect 21637 16739 21695 16745
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 24670 16736 24676 16788
rect 24728 16776 24734 16788
rect 24728 16748 25728 16776
rect 24728 16736 24734 16748
rect 25700 16708 25728 16748
rect 25774 16736 25780 16788
rect 25832 16776 25838 16788
rect 27433 16779 27491 16785
rect 27433 16776 27445 16779
rect 25832 16748 27445 16776
rect 25832 16736 25838 16748
rect 27433 16745 27445 16748
rect 27479 16745 27491 16779
rect 30098 16776 30104 16788
rect 27433 16739 27491 16745
rect 28460 16748 30104 16776
rect 21560 16680 22094 16708
rect 25700 16680 25820 16708
rect 17635 16612 18184 16640
rect 17635 16609 17647 16612
rect 17589 16603 17647 16609
rect 18230 16600 18236 16652
rect 18288 16640 18294 16652
rect 20806 16640 20812 16652
rect 18288 16612 18368 16640
rect 20767 16612 20812 16640
rect 18288 16600 18294 16612
rect 10873 16575 10931 16581
rect 10873 16541 10885 16575
rect 10919 16541 10931 16575
rect 10873 16535 10931 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 14921 16575 14979 16581
rect 14139 16544 14780 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 6420 16476 7604 16504
rect 10781 16507 10839 16513
rect 6420 16464 6426 16476
rect 10781 16473 10793 16507
rect 10827 16504 10839 16507
rect 10827 16476 11730 16504
rect 10827 16473 10839 16476
rect 10781 16467 10839 16473
rect 4525 16439 4583 16445
rect 4525 16405 4537 16439
rect 4571 16436 4583 16439
rect 4706 16436 4712 16448
rect 4571 16408 4712 16436
rect 4571 16405 4583 16408
rect 4525 16399 4583 16405
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 11330 16396 11336 16448
rect 11388 16436 11394 16448
rect 11425 16439 11483 16445
rect 11425 16436 11437 16439
rect 11388 16408 11437 16436
rect 11388 16396 11394 16408
rect 11425 16405 11437 16408
rect 11471 16405 11483 16439
rect 14274 16436 14280 16448
rect 14235 16408 14280 16436
rect 11425 16399 11483 16405
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 14752 16436 14780 16544
rect 14921 16541 14933 16575
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15381 16575 15439 16581
rect 15381 16541 15393 16575
rect 15427 16541 15439 16575
rect 15381 16535 15439 16541
rect 17862 16532 17868 16584
rect 17920 16572 17926 16584
rect 18340 16581 18368 16612
rect 20806 16600 20812 16612
rect 20864 16600 20870 16652
rect 21082 16640 21088 16652
rect 21043 16612 21088 16640
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21174 16600 21180 16652
rect 21232 16640 21238 16652
rect 22066 16640 22094 16680
rect 24397 16643 24455 16649
rect 24397 16640 24409 16643
rect 21232 16612 21956 16640
rect 22066 16612 24409 16640
rect 21232 16600 21238 16612
rect 18325 16575 18383 16581
rect 17920 16544 17965 16572
rect 17920 16532 17926 16544
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 21928 16572 21956 16612
rect 24397 16609 24409 16612
rect 24443 16609 24455 16643
rect 24397 16603 24455 16609
rect 24673 16643 24731 16649
rect 24673 16609 24685 16643
rect 24719 16640 24731 16643
rect 25406 16640 25412 16652
rect 24719 16612 25412 16640
rect 24719 16609 24731 16612
rect 24673 16603 24731 16609
rect 25406 16600 25412 16612
rect 25464 16600 25470 16652
rect 25792 16640 25820 16680
rect 25958 16668 25964 16720
rect 26016 16708 26022 16720
rect 28460 16717 28488 16748
rect 30098 16736 30104 16748
rect 30156 16736 30162 16788
rect 32769 16779 32827 16785
rect 31128 16748 32720 16776
rect 28445 16711 28503 16717
rect 28445 16708 28457 16711
rect 26016 16680 28457 16708
rect 26016 16668 26022 16680
rect 28445 16677 28457 16680
rect 28491 16677 28503 16711
rect 28445 16671 28503 16677
rect 28997 16711 29055 16717
rect 28997 16677 29009 16711
rect 29043 16708 29055 16711
rect 29043 16680 30052 16708
rect 29043 16677 29055 16680
rect 28997 16671 29055 16677
rect 29546 16640 29552 16652
rect 25792 16612 26648 16640
rect 29507 16612 29552 16640
rect 22097 16575 22155 16581
rect 22097 16572 22109 16575
rect 18472 16544 18517 16572
rect 21928 16544 22109 16572
rect 18472 16532 18478 16544
rect 22097 16541 22109 16544
rect 22143 16541 22155 16575
rect 22097 16535 22155 16541
rect 23474 16532 23480 16584
rect 23532 16532 23538 16584
rect 26620 16581 26648 16612
rect 29546 16600 29552 16612
rect 29604 16600 29610 16652
rect 30024 16649 30052 16680
rect 30009 16643 30067 16649
rect 30009 16609 30021 16643
rect 30055 16640 30067 16643
rect 31128 16640 31156 16748
rect 32692 16708 32720 16748
rect 32769 16745 32781 16779
rect 32815 16776 32827 16779
rect 33134 16776 33140 16788
rect 32815 16748 33140 16776
rect 32815 16745 32827 16748
rect 32769 16739 32827 16745
rect 33134 16736 33140 16748
rect 33192 16736 33198 16788
rect 33318 16776 33324 16788
rect 33279 16748 33324 16776
rect 33318 16736 33324 16748
rect 33376 16736 33382 16788
rect 35894 16736 35900 16788
rect 35952 16776 35958 16788
rect 39209 16779 39267 16785
rect 39209 16776 39221 16779
rect 35952 16748 39221 16776
rect 35952 16736 35958 16748
rect 39209 16745 39221 16748
rect 39255 16745 39267 16779
rect 39209 16739 39267 16745
rect 39758 16736 39764 16788
rect 39816 16776 39822 16788
rect 39945 16779 40003 16785
rect 39945 16776 39957 16779
rect 39816 16748 39957 16776
rect 39816 16736 39822 16748
rect 39945 16745 39957 16748
rect 39991 16745 40003 16779
rect 39945 16739 40003 16745
rect 40681 16779 40739 16785
rect 40681 16745 40693 16779
rect 40727 16776 40739 16779
rect 40770 16776 40776 16788
rect 40727 16748 40776 16776
rect 40727 16745 40739 16748
rect 40681 16739 40739 16745
rect 40770 16736 40776 16748
rect 40828 16736 40834 16788
rect 42794 16736 42800 16788
rect 42852 16776 42858 16788
rect 44082 16776 44088 16788
rect 42852 16748 44088 16776
rect 42852 16736 42858 16748
rect 44082 16736 44088 16748
rect 44140 16736 44146 16788
rect 44266 16736 44272 16788
rect 44324 16776 44330 16788
rect 47026 16776 47032 16788
rect 44324 16748 47032 16776
rect 44324 16736 44330 16748
rect 47026 16736 47032 16748
rect 47084 16776 47090 16788
rect 47121 16779 47179 16785
rect 47121 16776 47133 16779
rect 47084 16748 47133 16776
rect 47084 16736 47090 16748
rect 47121 16745 47133 16748
rect 47167 16745 47179 16779
rect 47121 16739 47179 16745
rect 35802 16708 35808 16720
rect 32692 16680 35808 16708
rect 35802 16668 35808 16680
rect 35860 16668 35866 16720
rect 31294 16640 31300 16652
rect 30055 16612 31156 16640
rect 31255 16612 31300 16640
rect 30055 16609 30067 16612
rect 30009 16603 30067 16609
rect 31294 16600 31300 16612
rect 31352 16600 31358 16652
rect 33962 16600 33968 16652
rect 34020 16640 34026 16652
rect 35912 16640 35940 16736
rect 41782 16668 41788 16720
rect 41840 16708 41846 16720
rect 43162 16708 43168 16720
rect 41840 16680 43168 16708
rect 41840 16668 41846 16680
rect 43162 16668 43168 16680
rect 43220 16668 43226 16720
rect 44910 16708 44916 16720
rect 43272 16680 44916 16708
rect 36354 16640 36360 16652
rect 34020 16612 35940 16640
rect 36315 16612 36360 16640
rect 34020 16600 34026 16612
rect 26605 16575 26663 16581
rect 26605 16541 26617 16575
rect 26651 16574 26663 16575
rect 27525 16575 27583 16581
rect 26651 16546 26685 16574
rect 26651 16541 26663 16546
rect 26605 16535 26663 16541
rect 27525 16541 27537 16575
rect 27571 16572 27583 16575
rect 27706 16572 27712 16584
rect 27571 16544 27712 16572
rect 27571 16541 27583 16544
rect 27525 16535 27583 16541
rect 27706 16532 27712 16544
rect 27764 16532 27770 16584
rect 28166 16532 28172 16584
rect 28224 16572 28230 16584
rect 28721 16575 28779 16581
rect 28721 16572 28733 16575
rect 28224 16544 28733 16572
rect 28224 16532 28230 16544
rect 28721 16541 28733 16544
rect 28767 16541 28779 16575
rect 28721 16535 28779 16541
rect 29730 16532 29736 16584
rect 29788 16572 29794 16584
rect 29917 16575 29975 16581
rect 29917 16572 29929 16575
rect 29788 16544 29929 16572
rect 29788 16532 29794 16544
rect 29917 16541 29929 16544
rect 29963 16541 29975 16575
rect 31018 16572 31024 16584
rect 30979 16544 31024 16572
rect 29917 16535 29975 16541
rect 14829 16507 14887 16513
rect 14829 16473 14841 16507
rect 14875 16504 14887 16507
rect 14875 16476 16422 16504
rect 14875 16473 14887 16476
rect 14829 16467 14887 16473
rect 18598 16464 18604 16516
rect 18656 16504 18662 16516
rect 18656 16476 19642 16504
rect 18656 16464 18662 16476
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 22373 16507 22431 16513
rect 22373 16504 22385 16507
rect 22336 16476 22385 16504
rect 22336 16464 22342 16476
rect 22373 16473 22385 16476
rect 22419 16473 22431 16507
rect 26697 16507 26755 16513
rect 26697 16504 26709 16507
rect 25898 16476 26709 16504
rect 22373 16467 22431 16473
rect 26697 16473 26709 16476
rect 26743 16473 26755 16507
rect 26697 16467 26755 16473
rect 15194 16436 15200 16448
rect 14752 16408 15200 16436
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 15473 16439 15531 16445
rect 15473 16405 15485 16439
rect 15519 16436 15531 16439
rect 15746 16436 15752 16448
rect 15519 16408 15752 16436
rect 15519 16405 15531 16408
rect 15473 16399 15531 16405
rect 15746 16396 15752 16408
rect 15804 16396 15810 16448
rect 16114 16436 16120 16448
rect 16075 16408 16120 16436
rect 16114 16396 16120 16408
rect 16172 16396 16178 16448
rect 16298 16396 16304 16448
rect 16356 16436 16362 16448
rect 19337 16439 19395 16445
rect 19337 16436 19349 16439
rect 16356 16408 19349 16436
rect 16356 16396 16362 16408
rect 19337 16405 19349 16408
rect 19383 16405 19395 16439
rect 19337 16399 19395 16405
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 23845 16439 23903 16445
rect 23845 16436 23857 16439
rect 21048 16408 23857 16436
rect 21048 16396 21054 16408
rect 23845 16405 23857 16408
rect 23891 16436 23903 16439
rect 24670 16436 24676 16448
rect 23891 16408 24676 16436
rect 23891 16405 23903 16408
rect 23845 16399 23903 16405
rect 24670 16396 24676 16408
rect 24728 16396 24734 16448
rect 26145 16439 26203 16445
rect 26145 16405 26157 16439
rect 26191 16436 26203 16439
rect 27614 16436 27620 16448
rect 26191 16408 27620 16436
rect 26191 16405 26203 16408
rect 26145 16399 26203 16405
rect 27614 16396 27620 16408
rect 27672 16396 27678 16448
rect 28626 16436 28632 16448
rect 28587 16408 28632 16436
rect 28626 16396 28632 16408
rect 28684 16396 28690 16448
rect 28810 16436 28816 16448
rect 28771 16408 28816 16436
rect 28810 16396 28816 16408
rect 28868 16396 28874 16448
rect 29932 16436 29960 16535
rect 31018 16532 31024 16544
rect 31076 16532 31082 16584
rect 34164 16581 34192 16612
rect 36354 16600 36360 16612
rect 36412 16600 36418 16652
rect 36633 16643 36691 16649
rect 36633 16609 36645 16643
rect 36679 16640 36691 16643
rect 37642 16640 37648 16652
rect 36679 16612 37648 16640
rect 36679 16609 36691 16612
rect 36633 16603 36691 16609
rect 37642 16600 37648 16612
rect 37700 16600 37706 16652
rect 38286 16600 38292 16652
rect 38344 16640 38350 16652
rect 38344 16612 38608 16640
rect 38344 16600 38350 16612
rect 34149 16575 34207 16581
rect 34149 16541 34161 16575
rect 34195 16541 34207 16575
rect 34790 16572 34796 16584
rect 34751 16544 34796 16572
rect 34149 16535 34207 16541
rect 34790 16532 34796 16544
rect 34848 16532 34854 16584
rect 34885 16575 34943 16581
rect 34885 16541 34897 16575
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 31754 16464 31760 16516
rect 31812 16464 31818 16516
rect 33413 16507 33471 16513
rect 33413 16473 33425 16507
rect 33459 16504 33471 16507
rect 34238 16504 34244 16516
rect 33459 16476 34244 16504
rect 33459 16473 33471 16476
rect 33413 16467 33471 16473
rect 34238 16464 34244 16476
rect 34296 16464 34302 16516
rect 34900 16504 34928 16535
rect 35342 16532 35348 16584
rect 35400 16572 35406 16584
rect 35437 16575 35495 16581
rect 35437 16572 35449 16575
rect 35400 16544 35449 16572
rect 35400 16532 35406 16544
rect 35437 16541 35449 16544
rect 35483 16541 35495 16575
rect 35437 16535 35495 16541
rect 35526 16532 35532 16584
rect 35584 16572 35590 16584
rect 38580 16581 38608 16612
rect 40678 16600 40684 16652
rect 40736 16640 40742 16652
rect 42610 16640 42616 16652
rect 40736 16612 40816 16640
rect 42571 16612 42616 16640
rect 40736 16600 40742 16612
rect 40788 16581 40816 16612
rect 42610 16600 42616 16612
rect 42668 16600 42674 16652
rect 43272 16581 43300 16680
rect 44910 16668 44916 16680
rect 44968 16668 44974 16720
rect 44174 16600 44180 16652
rect 44232 16640 44238 16652
rect 44232 16612 44588 16640
rect 44232 16600 44238 16612
rect 38565 16575 38623 16581
rect 35584 16544 35629 16572
rect 35584 16532 35590 16544
rect 38565 16541 38577 16575
rect 38611 16541 38623 16575
rect 38565 16535 38623 16541
rect 40037 16575 40095 16581
rect 40037 16541 40049 16575
rect 40083 16541 40095 16575
rect 40037 16535 40095 16541
rect 40773 16575 40831 16581
rect 40773 16541 40785 16575
rect 40819 16541 40831 16575
rect 40773 16535 40831 16541
rect 43257 16575 43315 16581
rect 43257 16541 43269 16575
rect 43303 16541 43315 16575
rect 43257 16535 43315 16541
rect 43717 16575 43775 16581
rect 43717 16541 43729 16575
rect 43763 16541 43775 16575
rect 44560 16572 44588 16612
rect 44634 16600 44640 16652
rect 44692 16640 44698 16652
rect 45649 16643 45707 16649
rect 45649 16640 45661 16643
rect 44692 16612 45661 16640
rect 44692 16600 44698 16612
rect 45649 16609 45661 16612
rect 45695 16609 45707 16643
rect 45649 16603 45707 16609
rect 45373 16575 45431 16581
rect 45373 16572 45385 16575
rect 44560 16544 45385 16572
rect 43717 16535 43775 16541
rect 45373 16541 45385 16544
rect 45419 16541 45431 16575
rect 45373 16535 45431 16541
rect 35544 16504 35572 16532
rect 38657 16507 38715 16513
rect 38657 16504 38669 16507
rect 34900 16476 35572 16504
rect 37858 16476 38669 16504
rect 38657 16473 38669 16476
rect 38703 16473 38715 16507
rect 38657 16467 38715 16473
rect 33870 16436 33876 16448
rect 29932 16408 33876 16436
rect 33870 16396 33876 16408
rect 33928 16396 33934 16448
rect 34054 16436 34060 16448
rect 34015 16408 34060 16436
rect 34054 16396 34060 16408
rect 34112 16396 34118 16448
rect 38105 16439 38163 16445
rect 38105 16405 38117 16439
rect 38151 16436 38163 16439
rect 40052 16436 40080 16535
rect 41506 16464 41512 16516
rect 41564 16504 41570 16516
rect 43073 16507 43131 16513
rect 43073 16504 43085 16507
rect 41564 16476 43085 16504
rect 41564 16464 41570 16476
rect 43073 16473 43085 16476
rect 43119 16473 43131 16507
rect 43073 16467 43131 16473
rect 41046 16436 41052 16448
rect 38151 16408 41052 16436
rect 38151 16405 38163 16408
rect 38105 16399 38163 16405
rect 41046 16396 41052 16408
rect 41104 16396 41110 16448
rect 41322 16396 41328 16448
rect 41380 16436 41386 16448
rect 43732 16436 43760 16535
rect 44082 16464 44088 16516
rect 44140 16504 44146 16516
rect 47136 16504 47164 16739
rect 48406 16736 48412 16788
rect 48464 16776 48470 16788
rect 48501 16779 48559 16785
rect 48501 16776 48513 16779
rect 48464 16748 48513 16776
rect 48464 16736 48470 16748
rect 48501 16745 48513 16748
rect 48547 16745 48559 16779
rect 50154 16776 50160 16788
rect 50115 16748 50160 16776
rect 48501 16739 48559 16745
rect 50154 16736 50160 16748
rect 50212 16736 50218 16788
rect 52454 16736 52460 16788
rect 52512 16776 52518 16788
rect 54294 16776 54300 16788
rect 52512 16748 53880 16776
rect 54255 16748 54300 16776
rect 52512 16736 52518 16748
rect 49053 16711 49111 16717
rect 49053 16677 49065 16711
rect 49099 16677 49111 16711
rect 49053 16671 49111 16677
rect 47762 16600 47768 16652
rect 47820 16640 47826 16652
rect 49068 16640 49096 16671
rect 51350 16668 51356 16720
rect 51408 16708 51414 16720
rect 51408 16680 52776 16708
rect 51408 16668 51414 16680
rect 47820 16612 49096 16640
rect 47820 16600 47826 16612
rect 48056 16581 48084 16612
rect 49142 16600 49148 16652
rect 49200 16640 49206 16652
rect 49329 16643 49387 16649
rect 49329 16640 49341 16643
rect 49200 16612 49341 16640
rect 49200 16600 49206 16612
rect 49329 16609 49341 16612
rect 49375 16609 49387 16643
rect 50614 16640 50620 16652
rect 50575 16612 50620 16640
rect 49329 16603 49387 16609
rect 50614 16600 50620 16612
rect 50672 16600 50678 16652
rect 51442 16640 51448 16652
rect 51403 16612 51448 16640
rect 51442 16600 51448 16612
rect 51500 16600 51506 16652
rect 51721 16643 51779 16649
rect 51721 16609 51733 16643
rect 51767 16609 51779 16643
rect 52748 16640 52776 16680
rect 52822 16668 52828 16720
rect 52880 16708 52886 16720
rect 53285 16711 53343 16717
rect 53285 16708 53297 16711
rect 52880 16680 53297 16708
rect 52880 16668 52886 16680
rect 53285 16677 53297 16680
rect 53331 16708 53343 16711
rect 53374 16708 53380 16720
rect 53331 16680 53380 16708
rect 53331 16677 53343 16680
rect 53285 16671 53343 16677
rect 53374 16668 53380 16680
rect 53432 16668 53438 16720
rect 53852 16640 53880 16748
rect 54294 16736 54300 16748
rect 54352 16736 54358 16788
rect 54386 16640 54392 16652
rect 52748 16612 53328 16640
rect 51721 16603 51779 16609
rect 48041 16575 48099 16581
rect 48041 16541 48053 16575
rect 48087 16541 48099 16575
rect 48314 16572 48320 16584
rect 48275 16544 48320 16572
rect 48041 16535 48099 16541
rect 48314 16532 48320 16544
rect 48372 16532 48378 16584
rect 48961 16575 49019 16581
rect 48961 16541 48973 16575
rect 49007 16572 49019 16575
rect 49050 16572 49056 16584
rect 49007 16544 49056 16572
rect 49007 16541 49019 16544
rect 48961 16535 49019 16541
rect 49050 16532 49056 16544
rect 49108 16532 49114 16584
rect 50525 16575 50583 16581
rect 50525 16541 50537 16575
rect 50571 16572 50583 16575
rect 51736 16572 51764 16603
rect 53300 16584 53328 16612
rect 53852 16612 54392 16640
rect 51994 16572 52000 16584
rect 50571 16544 52000 16572
rect 50571 16541 50583 16544
rect 50525 16535 50583 16541
rect 51994 16532 52000 16544
rect 52052 16572 52058 16584
rect 52052 16566 52868 16572
rect 52052 16544 53144 16566
rect 52052 16532 52058 16544
rect 52840 16538 53144 16544
rect 44140 16476 46138 16504
rect 47136 16476 48314 16504
rect 44140 16464 44146 16476
rect 45848 16448 45876 16476
rect 48286 16448 48314 16476
rect 52454 16464 52460 16516
rect 52512 16504 52518 16516
rect 52512 16476 53052 16504
rect 52512 16464 52518 16476
rect 43898 16436 43904 16448
rect 41380 16408 43760 16436
rect 43859 16408 43904 16436
rect 41380 16396 41386 16408
rect 43898 16396 43904 16408
rect 43956 16396 43962 16448
rect 45830 16396 45836 16448
rect 45888 16396 45894 16448
rect 48130 16436 48136 16448
rect 48091 16408 48136 16436
rect 48130 16396 48136 16408
rect 48188 16396 48194 16448
rect 48222 16396 48228 16448
rect 48280 16436 48314 16448
rect 49053 16439 49111 16445
rect 49053 16436 49065 16439
rect 48280 16408 49065 16436
rect 48280 16396 48286 16408
rect 49053 16405 49065 16408
rect 49099 16405 49111 16439
rect 49053 16399 49111 16405
rect 49145 16439 49203 16445
rect 49145 16405 49157 16439
rect 49191 16436 49203 16439
rect 49234 16436 49240 16448
rect 49191 16408 49240 16436
rect 49191 16405 49203 16408
rect 49145 16399 49203 16405
rect 49234 16396 49240 16408
rect 49292 16396 49298 16448
rect 52730 16436 52736 16448
rect 52691 16408 52736 16436
rect 52730 16396 52736 16408
rect 52788 16396 52794 16448
rect 52822 16396 52828 16448
rect 52880 16436 52886 16448
rect 53024 16445 53052 16476
rect 53116 16445 53144 16538
rect 53282 16532 53288 16584
rect 53340 16532 53346 16584
rect 53852 16581 53880 16612
rect 54386 16600 54392 16612
rect 54444 16600 54450 16652
rect 55398 16640 55404 16652
rect 55359 16612 55404 16640
rect 55398 16600 55404 16612
rect 55456 16600 55462 16652
rect 56318 16600 56324 16652
rect 56376 16640 56382 16652
rect 56413 16643 56471 16649
rect 56413 16640 56425 16643
rect 56376 16612 56425 16640
rect 56376 16600 56382 16612
rect 56413 16609 56425 16612
rect 56459 16609 56471 16643
rect 56686 16640 56692 16652
rect 56647 16612 56692 16640
rect 56413 16603 56471 16609
rect 56686 16600 56692 16612
rect 56744 16600 56750 16652
rect 53837 16575 53895 16581
rect 53837 16541 53849 16575
rect 53883 16541 53895 16575
rect 53837 16535 53895 16541
rect 53926 16532 53932 16584
rect 53984 16572 53990 16584
rect 54113 16575 54171 16581
rect 53984 16544 54029 16572
rect 53984 16532 53990 16544
rect 54113 16541 54125 16575
rect 54159 16572 54171 16575
rect 55214 16572 55220 16584
rect 54159 16544 55220 16572
rect 54159 16541 54171 16544
rect 54113 16535 54171 16541
rect 55214 16532 55220 16544
rect 55272 16532 55278 16584
rect 55490 16572 55496 16584
rect 55451 16544 55496 16572
rect 55490 16532 55496 16544
rect 55548 16532 55554 16584
rect 53190 16464 53196 16516
rect 53248 16504 53254 16516
rect 55508 16504 55536 16532
rect 53248 16476 55536 16504
rect 53248 16464 53254 16476
rect 57422 16464 57428 16516
rect 57480 16464 57486 16516
rect 52917 16439 52975 16445
rect 52917 16436 52929 16439
rect 52880 16408 52929 16436
rect 52880 16396 52886 16408
rect 52917 16405 52929 16408
rect 52963 16405 52975 16439
rect 52917 16399 52975 16405
rect 53009 16439 53067 16445
rect 53009 16405 53021 16439
rect 53055 16405 53067 16439
rect 53009 16399 53067 16405
rect 53101 16439 53159 16445
rect 53101 16405 53113 16439
rect 53147 16436 53159 16439
rect 54110 16436 54116 16448
rect 53147 16408 54116 16436
rect 53147 16405 53159 16408
rect 53101 16399 53159 16405
rect 54110 16396 54116 16408
rect 54168 16396 54174 16448
rect 55861 16439 55919 16445
rect 55861 16405 55873 16439
rect 55907 16436 55919 16439
rect 56594 16436 56600 16448
rect 55907 16408 56600 16436
rect 55907 16405 55919 16408
rect 55861 16399 55919 16405
rect 56594 16396 56600 16408
rect 56652 16396 56658 16448
rect 56778 16396 56784 16448
rect 56836 16436 56842 16448
rect 58161 16439 58219 16445
rect 58161 16436 58173 16439
rect 56836 16408 58173 16436
rect 56836 16396 56842 16408
rect 58161 16405 58173 16408
rect 58207 16405 58219 16439
rect 58161 16399 58219 16405
rect 1104 16346 58880 16368
rect 1104 16294 15398 16346
rect 15450 16294 15462 16346
rect 15514 16294 15526 16346
rect 15578 16294 15590 16346
rect 15642 16294 15654 16346
rect 15706 16294 29846 16346
rect 29898 16294 29910 16346
rect 29962 16294 29974 16346
rect 30026 16294 30038 16346
rect 30090 16294 30102 16346
rect 30154 16294 44294 16346
rect 44346 16294 44358 16346
rect 44410 16294 44422 16346
rect 44474 16294 44486 16346
rect 44538 16294 44550 16346
rect 44602 16294 58880 16346
rect 1104 16272 58880 16294
rect 3418 16232 3424 16244
rect 3331 16204 3424 16232
rect 3418 16192 3424 16204
rect 3476 16232 3482 16244
rect 9858 16232 9864 16244
rect 3476 16204 9864 16232
rect 3476 16192 3482 16204
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 14274 16192 14280 16244
rect 14332 16232 14338 16244
rect 18966 16232 18972 16244
rect 14332 16204 18972 16232
rect 14332 16192 14338 16204
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 23106 16232 23112 16244
rect 20088 16204 22094 16232
rect 3326 16124 3332 16176
rect 3384 16164 3390 16176
rect 4525 16167 4583 16173
rect 4525 16164 4537 16167
rect 3384 16136 4537 16164
rect 3384 16124 3390 16136
rect 4525 16133 4537 16136
rect 4571 16133 4583 16167
rect 6730 16164 6736 16176
rect 4525 16127 4583 16133
rect 4632 16136 6736 16164
rect 3973 16099 4031 16105
rect 3973 16065 3985 16099
rect 4019 16096 4031 16099
rect 4062 16096 4068 16108
rect 4019 16068 4068 16096
rect 4019 16065 4031 16068
rect 3973 16059 4031 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 4632 16105 4660 16136
rect 6730 16124 6736 16136
rect 6788 16124 6794 16176
rect 9950 16124 9956 16176
rect 10008 16124 10014 16176
rect 12250 16164 12256 16176
rect 12211 16136 12256 16164
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 12710 16124 12716 16176
rect 12768 16124 12774 16176
rect 15746 16124 15752 16176
rect 15804 16164 15810 16176
rect 19702 16164 19708 16176
rect 15804 16136 17526 16164
rect 19663 16136 19708 16164
rect 15804 16124 15810 16136
rect 19702 16124 19708 16136
rect 19760 16124 19766 16176
rect 20088 16164 20116 16204
rect 20162 16164 20168 16176
rect 20088 16136 20168 16164
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 22066 16164 22094 16204
rect 22940 16204 23112 16232
rect 22189 16167 22247 16173
rect 22189 16164 22201 16167
rect 22066 16136 22201 16164
rect 22189 16133 22201 16136
rect 22235 16133 22247 16167
rect 22189 16127 22247 16133
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16065 4675 16099
rect 4617 16059 4675 16065
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 5316 16068 5457 16096
rect 5316 16056 5322 16068
rect 5445 16065 5457 16068
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16096 6423 16099
rect 7190 16096 7196 16108
rect 6411 16068 7196 16096
rect 6411 16065 6423 16068
rect 6365 16059 6423 16065
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 8757 16099 8815 16105
rect 8757 16065 8769 16099
rect 8803 16065 8815 16099
rect 14366 16096 14372 16108
rect 14327 16068 14372 16096
rect 8757 16059 8815 16065
rect 5350 16028 5356 16040
rect 5311 16000 5356 16028
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 8772 16028 8800 16059
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 22278 16056 22284 16108
rect 22336 16096 22342 16108
rect 22940 16105 22968 16204
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 29730 16232 29736 16244
rect 24596 16204 29736 16232
rect 23198 16164 23204 16176
rect 23159 16136 23204 16164
rect 23198 16124 23204 16136
rect 23256 16124 23262 16176
rect 24486 16164 24492 16176
rect 24426 16136 24492 16164
rect 24486 16124 24492 16136
rect 24544 16124 24550 16176
rect 22373 16099 22431 16105
rect 22373 16096 22385 16099
rect 22336 16068 22385 16096
rect 22336 16056 22342 16068
rect 22373 16065 22385 16068
rect 22419 16065 22431 16099
rect 22373 16059 22431 16065
rect 22925 16099 22983 16105
rect 22925 16065 22937 16099
rect 22971 16065 22983 16099
rect 22925 16059 22983 16065
rect 10594 16028 10600 16040
rect 8772 16000 10600 16028
rect 10594 15988 10600 16000
rect 10652 15988 10658 16040
rect 10686 15988 10692 16040
rect 10744 16028 10750 16040
rect 10965 16031 11023 16037
rect 10965 16028 10977 16031
rect 10744 16000 10977 16028
rect 10744 15988 10750 16000
rect 10965 15997 10977 16000
rect 11011 15997 11023 16031
rect 11974 16028 11980 16040
rect 11935 16000 11980 16028
rect 10965 15991 11023 15997
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 16298 16028 16304 16040
rect 13044 16000 16304 16028
rect 13044 15988 13050 16000
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 17218 16028 17224 16040
rect 17179 16000 17224 16028
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 18690 16028 18696 16040
rect 18651 16000 18696 16028
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 18969 16031 19027 16037
rect 18969 15997 18981 16031
rect 19015 15997 19027 16031
rect 19426 16028 19432 16040
rect 19387 16000 19432 16028
rect 18969 15991 19027 15997
rect 5810 15960 5816 15972
rect 5771 15932 5816 15960
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 6454 15960 6460 15972
rect 6415 15932 6460 15960
rect 6454 15920 6460 15932
rect 6512 15920 6518 15972
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 9217 15963 9275 15969
rect 9217 15960 9229 15963
rect 6788 15932 9229 15960
rect 6788 15920 6794 15932
rect 9217 15929 9229 15932
rect 9263 15929 9275 15963
rect 9217 15923 9275 15929
rect 13725 15963 13783 15969
rect 13725 15929 13737 15963
rect 13771 15960 13783 15963
rect 14734 15960 14740 15972
rect 13771 15932 14740 15960
rect 13771 15929 13783 15932
rect 13725 15923 13783 15929
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 18984 15960 19012 15991
rect 19426 15988 19432 16000
rect 19484 15988 19490 16040
rect 20254 16028 20260 16040
rect 19536 16000 20260 16028
rect 19536 15960 19564 16000
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 21177 16031 21235 16037
rect 21177 15997 21189 16031
rect 21223 16028 21235 16031
rect 24596 16028 24624 16204
rect 29730 16192 29736 16204
rect 29788 16192 29794 16244
rect 31481 16235 31539 16241
rect 31481 16201 31493 16235
rect 31527 16232 31539 16235
rect 31754 16232 31760 16244
rect 31527 16204 31760 16232
rect 31527 16201 31539 16204
rect 31481 16195 31539 16201
rect 31754 16192 31760 16204
rect 31812 16192 31818 16244
rect 33873 16235 33931 16241
rect 33873 16232 33885 16235
rect 32784 16204 33885 16232
rect 24670 16124 24676 16176
rect 24728 16164 24734 16176
rect 28074 16164 28080 16176
rect 24728 16136 28080 16164
rect 24728 16124 24734 16136
rect 28074 16124 28080 16136
rect 28132 16124 28138 16176
rect 32784 16164 32812 16204
rect 33873 16201 33885 16204
rect 33919 16201 33931 16235
rect 33873 16195 33931 16201
rect 37642 16192 37648 16244
rect 37700 16232 37706 16244
rect 37737 16235 37795 16241
rect 37737 16232 37749 16235
rect 37700 16204 37749 16232
rect 37700 16192 37706 16204
rect 37737 16201 37749 16204
rect 37783 16201 37795 16235
rect 39390 16232 39396 16244
rect 37737 16195 37795 16201
rect 38488 16204 39396 16232
rect 34054 16164 34060 16176
rect 30760 16136 32812 16164
rect 33626 16136 34060 16164
rect 25409 16099 25467 16105
rect 25409 16065 25421 16099
rect 25455 16096 25467 16099
rect 26602 16096 26608 16108
rect 25455 16068 26608 16096
rect 25455 16065 25467 16068
rect 25409 16059 25467 16065
rect 26602 16056 26608 16068
rect 26660 16056 26666 16108
rect 27614 16096 27620 16108
rect 27575 16068 27620 16096
rect 27614 16056 27620 16068
rect 27672 16056 27678 16108
rect 30760 16105 30788 16136
rect 34054 16124 34060 16136
rect 34112 16124 34118 16176
rect 34885 16167 34943 16173
rect 34885 16133 34897 16167
rect 34931 16164 34943 16167
rect 35250 16164 35256 16176
rect 34931 16136 35256 16164
rect 34931 16133 34943 16136
rect 34885 16127 34943 16133
rect 35250 16124 35256 16136
rect 35308 16124 35314 16176
rect 38488 16164 38516 16204
rect 39390 16192 39396 16204
rect 39448 16192 39454 16244
rect 41690 16192 41696 16244
rect 41748 16232 41754 16244
rect 45646 16232 45652 16244
rect 41748 16204 44036 16232
rect 41748 16192 41754 16204
rect 39117 16167 39175 16173
rect 39117 16164 39129 16167
rect 35452 16136 38516 16164
rect 38580 16136 39129 16164
rect 28997 16099 29055 16105
rect 28997 16096 29009 16099
rect 28000 16068 29009 16096
rect 27706 16028 27712 16040
rect 21223 16000 24624 16028
rect 27667 16000 27712 16028
rect 21223 15997 21235 16000
rect 21177 15991 21235 15997
rect 27706 15988 27712 16000
rect 27764 15988 27770 16040
rect 26053 15963 26111 15969
rect 26053 15960 26065 15963
rect 18984 15932 19564 15960
rect 24228 15932 26065 15960
rect 7469 15895 7527 15901
rect 7469 15861 7481 15895
rect 7515 15892 7527 15895
rect 7926 15892 7932 15904
rect 7515 15864 7932 15892
rect 7515 15861 7527 15864
rect 7469 15855 7527 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 10701 15895 10759 15901
rect 10701 15892 10713 15895
rect 8904 15864 10713 15892
rect 8904 15852 8910 15864
rect 10701 15861 10713 15864
rect 10747 15861 10759 15895
rect 10701 15855 10759 15861
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15344 15864 15669 15892
rect 15344 15852 15350 15864
rect 15657 15861 15669 15864
rect 15703 15861 15715 15895
rect 15657 15855 15715 15861
rect 16114 15852 16120 15904
rect 16172 15892 16178 15904
rect 20990 15892 20996 15904
rect 16172 15864 20996 15892
rect 16172 15852 16178 15864
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 21082 15852 21088 15904
rect 21140 15892 21146 15904
rect 24228 15892 24256 15932
rect 26053 15929 26065 15932
rect 26099 15960 26111 15963
rect 27338 15960 27344 15972
rect 26099 15932 27344 15960
rect 26099 15929 26111 15932
rect 26053 15923 26111 15929
rect 27338 15920 27344 15932
rect 27396 15920 27402 15972
rect 27522 15920 27528 15972
rect 27580 15960 27586 15972
rect 28000 15960 28028 16068
rect 28997 16065 29009 16068
rect 29043 16065 29055 16099
rect 28997 16059 29055 16065
rect 29365 16099 29423 16105
rect 29365 16065 29377 16099
rect 29411 16096 29423 16099
rect 30745 16099 30803 16105
rect 30745 16096 30757 16099
rect 29411 16068 30757 16096
rect 29411 16065 29423 16068
rect 29365 16059 29423 16065
rect 30745 16065 30757 16068
rect 30791 16065 30803 16099
rect 30745 16059 30803 16065
rect 30926 16056 30932 16108
rect 30984 16096 30990 16108
rect 31389 16099 31447 16105
rect 31389 16096 31401 16099
rect 30984 16068 31401 16096
rect 30984 16056 30990 16068
rect 31389 16065 31401 16068
rect 31435 16065 31447 16099
rect 31389 16059 31447 16065
rect 28445 16031 28503 16037
rect 28445 15997 28457 16031
rect 28491 16028 28503 16031
rect 29270 16028 29276 16040
rect 28491 16000 29276 16028
rect 28491 15997 28503 16000
rect 28445 15991 28503 15997
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 30009 16031 30067 16037
rect 30009 15997 30021 16031
rect 30055 16028 30067 16031
rect 30558 16028 30564 16040
rect 30055 16000 30564 16028
rect 30055 15997 30067 16000
rect 30009 15991 30067 15997
rect 30558 15988 30564 16000
rect 30616 15988 30622 16040
rect 32122 16028 32128 16040
rect 32083 16000 32128 16028
rect 32122 15988 32128 16000
rect 32180 15988 32186 16040
rect 32398 16028 32404 16040
rect 32359 16000 32404 16028
rect 32398 15988 32404 16000
rect 32456 15988 32462 16040
rect 33134 15988 33140 16040
rect 33192 16028 33198 16040
rect 35452 16028 35480 16136
rect 35989 16099 36047 16105
rect 35989 16065 36001 16099
rect 36035 16096 36047 16099
rect 36262 16096 36268 16108
rect 36035 16068 36268 16096
rect 36035 16065 36047 16068
rect 35989 16059 36047 16065
rect 36262 16056 36268 16068
rect 36320 16056 36326 16108
rect 38396 16105 38424 16136
rect 38580 16108 38608 16136
rect 39117 16133 39129 16136
rect 39163 16133 39175 16167
rect 39117 16127 39175 16133
rect 42058 16124 42064 16176
rect 42116 16164 42122 16176
rect 42116 16136 43194 16164
rect 42116 16124 42122 16136
rect 37829 16099 37887 16105
rect 37829 16065 37841 16099
rect 37875 16065 37887 16099
rect 37829 16059 37887 16065
rect 38381 16099 38439 16105
rect 38381 16065 38393 16099
rect 38427 16065 38439 16099
rect 38562 16096 38568 16108
rect 38523 16068 38568 16096
rect 38381 16059 38439 16065
rect 33192 16000 35480 16028
rect 33192 15988 33198 16000
rect 35802 15988 35808 16040
rect 35860 16028 35866 16040
rect 35897 16031 35955 16037
rect 35897 16028 35909 16031
rect 35860 16000 35909 16028
rect 35860 15988 35866 16000
rect 35897 15997 35909 16000
rect 35943 15997 35955 16031
rect 35897 15991 35955 15997
rect 36170 15988 36176 16040
rect 36228 16028 36234 16040
rect 36357 16031 36415 16037
rect 36357 16028 36369 16031
rect 36228 16000 36369 16028
rect 36228 15988 36234 16000
rect 36357 15997 36369 16000
rect 36403 15997 36415 16031
rect 37844 16028 37872 16059
rect 38562 16056 38568 16068
rect 38620 16056 38626 16108
rect 39022 16096 39028 16108
rect 38983 16068 39028 16096
rect 39022 16056 39028 16068
rect 39080 16056 39086 16108
rect 39666 16096 39672 16108
rect 39627 16068 39672 16096
rect 39666 16056 39672 16068
rect 39724 16056 39730 16108
rect 41046 16096 41052 16108
rect 41007 16068 41052 16096
rect 41046 16056 41052 16068
rect 41104 16056 41110 16108
rect 44008 16096 44036 16204
rect 44744 16204 45652 16232
rect 44744 16173 44772 16204
rect 45646 16192 45652 16204
rect 45704 16232 45710 16244
rect 46842 16232 46848 16244
rect 45704 16204 46848 16232
rect 45704 16192 45710 16204
rect 46842 16192 46848 16204
rect 46900 16192 46906 16244
rect 48130 16192 48136 16244
rect 48188 16232 48194 16244
rect 49237 16235 49295 16241
rect 49237 16232 49249 16235
rect 48188 16204 49249 16232
rect 48188 16192 48194 16204
rect 49237 16201 49249 16204
rect 49283 16201 49295 16235
rect 49237 16195 49295 16201
rect 50062 16192 50068 16244
rect 50120 16232 50126 16244
rect 50249 16235 50307 16241
rect 50249 16232 50261 16235
rect 50120 16204 50261 16232
rect 50120 16192 50126 16204
rect 50249 16201 50261 16204
rect 50295 16201 50307 16235
rect 50249 16195 50307 16201
rect 52454 16192 52460 16244
rect 52512 16232 52518 16244
rect 54202 16232 54208 16244
rect 52512 16204 54208 16232
rect 52512 16192 52518 16204
rect 54202 16192 54208 16204
rect 54260 16192 54266 16244
rect 55125 16235 55183 16241
rect 55125 16201 55137 16235
rect 55171 16232 55183 16235
rect 55398 16232 55404 16244
rect 55171 16204 55404 16232
rect 55171 16201 55183 16204
rect 55125 16195 55183 16201
rect 55398 16192 55404 16204
rect 55456 16192 55462 16244
rect 44729 16167 44787 16173
rect 44729 16133 44741 16167
rect 44775 16133 44787 16167
rect 44729 16127 44787 16133
rect 44945 16167 45003 16173
rect 44945 16133 44957 16167
rect 44991 16164 45003 16167
rect 45186 16164 45192 16176
rect 44991 16136 45192 16164
rect 44991 16133 45003 16136
rect 44945 16127 45003 16133
rect 45186 16124 45192 16136
rect 45244 16124 45250 16176
rect 45554 16164 45560 16176
rect 45515 16136 45560 16164
rect 45554 16124 45560 16136
rect 45612 16124 45618 16176
rect 48041 16167 48099 16173
rect 45664 16136 46796 16164
rect 45664 16096 45692 16136
rect 45830 16096 45836 16108
rect 44008 16068 45692 16096
rect 45791 16068 45836 16096
rect 45830 16056 45836 16068
rect 45888 16056 45894 16108
rect 46474 16096 46480 16108
rect 46435 16068 46480 16096
rect 46474 16056 46480 16068
rect 46532 16056 46538 16108
rect 46768 16040 46796 16136
rect 48041 16133 48053 16167
rect 48087 16164 48099 16167
rect 48958 16164 48964 16176
rect 48087 16136 48964 16164
rect 48087 16133 48099 16136
rect 48041 16127 48099 16133
rect 48958 16124 48964 16136
rect 49016 16124 49022 16176
rect 50893 16167 50951 16173
rect 50893 16133 50905 16167
rect 50939 16164 50951 16167
rect 51813 16167 51871 16173
rect 51813 16164 51825 16167
rect 50939 16136 51825 16164
rect 50939 16133 50951 16136
rect 50893 16127 50951 16133
rect 51813 16133 51825 16136
rect 51859 16164 51871 16167
rect 51859 16136 52868 16164
rect 51859 16133 51871 16136
rect 51813 16127 51871 16133
rect 47949 16099 48007 16105
rect 47949 16065 47961 16099
rect 47995 16065 48007 16099
rect 47949 16059 48007 16065
rect 40957 16031 41015 16037
rect 40957 16028 40969 16031
rect 37844 16000 40969 16028
rect 36357 15991 36415 15997
rect 40957 15997 40969 16000
rect 41003 16028 41015 16031
rect 41230 16028 41236 16040
rect 41003 16000 41236 16028
rect 41003 15997 41015 16000
rect 40957 15991 41015 15997
rect 41230 15988 41236 16000
rect 41288 15988 41294 16040
rect 41874 16028 41880 16040
rect 41835 16000 41880 16028
rect 41874 15988 41880 16000
rect 41932 15988 41938 16040
rect 42429 16031 42487 16037
rect 42429 15997 42441 16031
rect 42475 15997 42487 16031
rect 42429 15991 42487 15997
rect 42705 16031 42763 16037
rect 42705 15997 42717 16031
rect 42751 16028 42763 16031
rect 44174 16028 44180 16040
rect 42751 16000 44180 16028
rect 42751 15997 42763 16000
rect 42705 15991 42763 15997
rect 27580 15932 28028 15960
rect 27580 15920 27586 15932
rect 33870 15920 33876 15972
rect 33928 15960 33934 15972
rect 38838 15960 38844 15972
rect 33928 15932 38844 15960
rect 33928 15920 33934 15932
rect 38838 15920 38844 15932
rect 38896 15920 38902 15972
rect 39022 15920 39028 15972
rect 39080 15960 39086 15972
rect 39761 15963 39819 15969
rect 39761 15960 39773 15963
rect 39080 15932 39773 15960
rect 39080 15920 39086 15932
rect 39761 15929 39773 15932
rect 39807 15960 39819 15963
rect 42444 15960 42472 15991
rect 44174 15988 44180 16000
rect 44232 15988 44238 16040
rect 46750 15988 46756 16040
rect 46808 16028 46814 16040
rect 47964 16028 47992 16059
rect 48130 16056 48136 16108
rect 48188 16096 48194 16108
rect 48225 16099 48283 16105
rect 48225 16096 48237 16099
rect 48188 16068 48237 16096
rect 48188 16056 48194 16068
rect 48225 16065 48237 16068
rect 48271 16096 48283 16099
rect 48314 16096 48320 16108
rect 48271 16068 48320 16096
rect 48271 16065 48283 16068
rect 48225 16059 48283 16065
rect 48314 16056 48320 16068
rect 48372 16056 48378 16108
rect 48869 16099 48927 16105
rect 48869 16065 48881 16099
rect 48915 16065 48927 16099
rect 48869 16059 48927 16065
rect 49053 16099 49111 16105
rect 49053 16065 49065 16099
rect 49099 16096 49111 16099
rect 49326 16096 49332 16108
rect 49099 16068 49332 16096
rect 49099 16065 49111 16068
rect 49053 16059 49111 16065
rect 48038 16028 48044 16040
rect 46808 16000 46853 16028
rect 47964 16000 48044 16028
rect 46808 15988 46814 16000
rect 48038 15988 48044 16000
rect 48096 16028 48102 16040
rect 48884 16028 48912 16059
rect 49326 16056 49332 16068
rect 49384 16056 49390 16108
rect 50985 16099 51043 16105
rect 50985 16065 50997 16099
rect 51031 16096 51043 16099
rect 51350 16096 51356 16108
rect 51031 16068 51356 16096
rect 51031 16065 51043 16068
rect 50985 16059 51043 16065
rect 51350 16056 51356 16068
rect 51408 16056 51414 16108
rect 51905 16099 51963 16105
rect 51905 16065 51917 16099
rect 51951 16096 51963 16099
rect 52730 16096 52736 16108
rect 51951 16068 52736 16096
rect 51951 16065 51963 16068
rect 51905 16059 51963 16065
rect 52730 16056 52736 16068
rect 52788 16056 52794 16108
rect 52840 16105 52868 16136
rect 53374 16124 53380 16176
rect 53432 16164 53438 16176
rect 53558 16164 53564 16176
rect 53432 16136 53564 16164
rect 53432 16124 53438 16136
rect 53558 16124 53564 16136
rect 53616 16164 53622 16176
rect 53837 16167 53895 16173
rect 53837 16164 53849 16167
rect 53616 16136 53849 16164
rect 53616 16124 53622 16136
rect 53837 16133 53849 16136
rect 53883 16133 53895 16167
rect 55953 16167 56011 16173
rect 55953 16164 55965 16167
rect 53837 16127 53895 16133
rect 54680 16136 55965 16164
rect 52825 16099 52883 16105
rect 52825 16065 52837 16099
rect 52871 16065 52883 16099
rect 52825 16059 52883 16065
rect 53653 16099 53711 16105
rect 53653 16065 53665 16099
rect 53699 16096 53711 16099
rect 54110 16096 54116 16108
rect 53699 16068 54116 16096
rect 53699 16065 53711 16068
rect 53653 16059 53711 16065
rect 54110 16056 54116 16068
rect 54168 16056 54174 16108
rect 54680 16105 54708 16136
rect 55953 16133 55965 16136
rect 55999 16133 56011 16167
rect 55953 16127 56011 16133
rect 54665 16099 54723 16105
rect 54665 16065 54677 16099
rect 54711 16065 54723 16099
rect 54665 16059 54723 16065
rect 54754 16056 54760 16108
rect 54812 16096 54818 16108
rect 54812 16068 54857 16096
rect 54812 16056 54818 16068
rect 54938 16056 54944 16108
rect 54996 16096 55002 16108
rect 55585 16099 55643 16105
rect 54996 16068 55041 16096
rect 54996 16056 55002 16068
rect 55585 16065 55597 16099
rect 55631 16065 55643 16099
rect 55585 16059 55643 16065
rect 48096 16000 48912 16028
rect 52089 16031 52147 16037
rect 48096 15988 48102 16000
rect 52089 15997 52101 16031
rect 52135 15997 52147 16031
rect 52089 15991 52147 15997
rect 46014 15960 46020 15972
rect 39807 15932 42472 15960
rect 45020 15932 46020 15960
rect 39807 15929 39819 15932
rect 39761 15923 39819 15929
rect 45020 15904 45048 15932
rect 46014 15920 46020 15932
rect 46072 15920 46078 15972
rect 48222 15920 48228 15972
rect 48280 15960 48286 15972
rect 52104 15960 52132 15991
rect 52546 15988 52552 16040
rect 52604 16028 52610 16040
rect 53009 16031 53067 16037
rect 53009 16028 53021 16031
rect 52604 16000 53021 16028
rect 52604 15988 52610 16000
rect 53009 15997 53021 16000
rect 53055 15997 53067 16031
rect 53009 15991 53067 15997
rect 54021 16031 54079 16037
rect 54021 15997 54033 16031
rect 54067 16028 54079 16031
rect 55030 16028 55036 16040
rect 54067 16000 55036 16028
rect 54067 15997 54079 16000
rect 54021 15991 54079 15997
rect 55030 15988 55036 16000
rect 55088 16028 55094 16040
rect 55600 16028 55628 16059
rect 55766 16056 55772 16108
rect 55824 16096 55830 16108
rect 56410 16096 56416 16108
rect 55824 16068 56416 16096
rect 55824 16056 55830 16068
rect 56410 16056 56416 16068
rect 56468 16056 56474 16108
rect 57146 16096 57152 16108
rect 57107 16068 57152 16096
rect 57146 16056 57152 16068
rect 57204 16056 57210 16108
rect 57054 16028 57060 16040
rect 55088 16000 55628 16028
rect 57015 16000 57060 16028
rect 55088 15988 55094 16000
rect 57054 15988 57060 16000
rect 57112 15988 57118 16040
rect 53190 15960 53196 15972
rect 48280 15932 48912 15960
rect 52104 15932 53196 15960
rect 48280 15920 48286 15932
rect 21140 15864 24256 15892
rect 21140 15852 21146 15864
rect 24394 15852 24400 15904
rect 24452 15892 24458 15904
rect 24673 15895 24731 15901
rect 24673 15892 24685 15895
rect 24452 15864 24685 15892
rect 24452 15852 24458 15864
rect 24673 15861 24685 15864
rect 24719 15861 24731 15895
rect 24673 15855 24731 15861
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 25501 15895 25559 15901
rect 25501 15892 25513 15895
rect 25464 15864 25513 15892
rect 25464 15852 25470 15864
rect 25501 15861 25513 15864
rect 25547 15861 25559 15895
rect 25501 15855 25559 15861
rect 30374 15852 30380 15904
rect 30432 15892 30438 15904
rect 30653 15895 30711 15901
rect 30653 15892 30665 15895
rect 30432 15864 30665 15892
rect 30432 15852 30438 15864
rect 30653 15861 30665 15864
rect 30699 15861 30711 15895
rect 30653 15855 30711 15861
rect 34882 15852 34888 15904
rect 34940 15892 34946 15904
rect 34977 15895 35035 15901
rect 34977 15892 34989 15895
rect 34940 15864 34989 15892
rect 34940 15852 34946 15864
rect 34977 15861 34989 15864
rect 35023 15861 35035 15895
rect 38562 15892 38568 15904
rect 38523 15864 38568 15892
rect 34977 15855 35035 15861
rect 38562 15852 38568 15864
rect 38620 15852 38626 15904
rect 44177 15895 44235 15901
rect 44177 15861 44189 15895
rect 44223 15892 44235 15895
rect 44726 15892 44732 15904
rect 44223 15864 44732 15892
rect 44223 15861 44235 15864
rect 44177 15855 44235 15861
rect 44726 15852 44732 15864
rect 44784 15852 44790 15904
rect 44913 15895 44971 15901
rect 44913 15861 44925 15895
rect 44959 15892 44971 15895
rect 45002 15892 45008 15904
rect 44959 15864 45008 15892
rect 44959 15861 44971 15864
rect 44913 15855 44971 15861
rect 45002 15852 45008 15864
rect 45060 15852 45066 15904
rect 45097 15895 45155 15901
rect 45097 15861 45109 15895
rect 45143 15892 45155 15895
rect 45554 15892 45560 15904
rect 45143 15864 45560 15892
rect 45143 15861 45155 15864
rect 45097 15855 45155 15861
rect 45554 15852 45560 15864
rect 45612 15852 45618 15904
rect 48314 15852 48320 15904
rect 48372 15892 48378 15904
rect 48884 15901 48912 15932
rect 53190 15920 53196 15932
rect 53248 15920 53254 15972
rect 56686 15920 56692 15972
rect 56744 15960 56750 15972
rect 56781 15963 56839 15969
rect 56781 15960 56793 15963
rect 56744 15932 56793 15960
rect 56744 15920 56750 15932
rect 56781 15929 56793 15932
rect 56827 15929 56839 15963
rect 56781 15923 56839 15929
rect 48409 15895 48467 15901
rect 48409 15892 48421 15895
rect 48372 15864 48421 15892
rect 48372 15852 48378 15864
rect 48409 15861 48421 15864
rect 48455 15861 48467 15895
rect 48409 15855 48467 15861
rect 48869 15895 48927 15901
rect 48869 15861 48881 15895
rect 48915 15861 48927 15895
rect 49694 15892 49700 15904
rect 49655 15864 49700 15892
rect 48869 15855 48927 15861
rect 49694 15852 49700 15864
rect 49752 15852 49758 15904
rect 51258 15852 51264 15904
rect 51316 15892 51322 15904
rect 51445 15895 51503 15901
rect 51445 15892 51457 15895
rect 51316 15864 51457 15892
rect 51316 15852 51322 15864
rect 51445 15861 51457 15864
rect 51491 15861 51503 15895
rect 51445 15855 51503 15861
rect 52917 15895 52975 15901
rect 52917 15861 52929 15895
rect 52963 15892 52975 15895
rect 53742 15892 53748 15904
rect 52963 15864 53748 15892
rect 52963 15861 52975 15864
rect 52917 15855 52975 15861
rect 53742 15852 53748 15864
rect 53800 15852 53806 15904
rect 1104 15802 58880 15824
rect 1104 15750 8174 15802
rect 8226 15750 8238 15802
rect 8290 15750 8302 15802
rect 8354 15750 8366 15802
rect 8418 15750 8430 15802
rect 8482 15750 22622 15802
rect 22674 15750 22686 15802
rect 22738 15750 22750 15802
rect 22802 15750 22814 15802
rect 22866 15750 22878 15802
rect 22930 15750 37070 15802
rect 37122 15750 37134 15802
rect 37186 15750 37198 15802
rect 37250 15750 37262 15802
rect 37314 15750 37326 15802
rect 37378 15750 51518 15802
rect 51570 15750 51582 15802
rect 51634 15750 51646 15802
rect 51698 15750 51710 15802
rect 51762 15750 51774 15802
rect 51826 15750 58880 15802
rect 1104 15728 58880 15750
rect 9122 15688 9128 15700
rect 9083 15660 9128 15688
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 10962 15688 10968 15700
rect 10652 15660 10968 15688
rect 10652 15648 10658 15660
rect 10962 15648 10968 15660
rect 11020 15688 11026 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 11020 15660 12357 15688
rect 11020 15648 11026 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 12345 15651 12403 15657
rect 14645 15691 14703 15697
rect 14645 15657 14657 15691
rect 14691 15688 14703 15691
rect 16482 15688 16488 15700
rect 14691 15660 16488 15688
rect 14691 15657 14703 15660
rect 14645 15651 14703 15657
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 18598 15688 18604 15700
rect 18559 15660 18604 15688
rect 18598 15648 18604 15660
rect 18656 15648 18662 15700
rect 19337 15691 19395 15697
rect 19337 15657 19349 15691
rect 19383 15688 19395 15691
rect 20622 15688 20628 15700
rect 19383 15660 20628 15688
rect 19383 15657 19395 15660
rect 19337 15651 19395 15657
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 23842 15688 23848 15700
rect 23803 15660 23848 15688
rect 23842 15648 23848 15660
rect 23900 15648 23906 15700
rect 24486 15688 24492 15700
rect 24447 15660 24492 15688
rect 24486 15648 24492 15660
rect 24544 15648 24550 15700
rect 26234 15688 26240 15700
rect 24596 15660 26240 15688
rect 5626 15580 5632 15632
rect 5684 15620 5690 15632
rect 9769 15623 9827 15629
rect 5684 15592 9444 15620
rect 5684 15580 5690 15592
rect 6178 15512 6184 15564
rect 6236 15552 6242 15564
rect 8294 15552 8300 15564
rect 6236 15524 6776 15552
rect 8255 15524 8300 15552
rect 6236 15512 6242 15524
rect 6748 15496 6776 15524
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 8754 15512 8760 15564
rect 8812 15552 8818 15564
rect 8812 15524 9260 15552
rect 8812 15512 8818 15524
rect 9232 15496 9260 15524
rect 5353 15487 5411 15493
rect 5353 15453 5365 15487
rect 5399 15453 5411 15487
rect 5353 15447 5411 15453
rect 5368 15416 5396 15447
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 5500 15456 5545 15484
rect 5500 15444 5506 15456
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 6546 15484 6552 15496
rect 6144 15456 6552 15484
rect 6144 15444 6150 15456
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 8389 15487 8447 15493
rect 6788 15456 6881 15484
rect 6788 15444 6794 15456
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 9122 15484 9128 15496
rect 8435 15456 9128 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 9416 15484 9444 15592
rect 9769 15589 9781 15623
rect 9815 15620 9827 15623
rect 11054 15620 11060 15632
rect 9815 15592 11060 15620
rect 9815 15589 9827 15592
rect 9769 15583 9827 15589
rect 11054 15580 11060 15592
rect 11112 15580 11118 15632
rect 15197 15623 15255 15629
rect 15197 15589 15209 15623
rect 15243 15589 15255 15623
rect 15197 15583 15255 15589
rect 17957 15623 18015 15629
rect 17957 15589 17969 15623
rect 18003 15620 18015 15623
rect 19426 15620 19432 15632
rect 18003 15592 19432 15620
rect 18003 15589 18015 15592
rect 17957 15583 18015 15589
rect 9490 15512 9496 15564
rect 9548 15552 9554 15564
rect 12986 15552 12992 15564
rect 9548 15524 12992 15552
rect 9548 15512 9554 15524
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 15212 15552 15240 15583
rect 19426 15580 19432 15592
rect 19484 15580 19490 15632
rect 24596 15620 24624 15660
rect 26234 15648 26240 15660
rect 26292 15648 26298 15700
rect 28261 15691 28319 15697
rect 28261 15657 28273 15691
rect 28307 15688 28319 15691
rect 32398 15688 32404 15700
rect 28307 15660 32404 15688
rect 28307 15657 28319 15660
rect 28261 15651 28319 15657
rect 32398 15648 32404 15660
rect 32456 15648 32462 15700
rect 36354 15648 36360 15700
rect 36412 15688 36418 15700
rect 36449 15691 36507 15697
rect 36449 15688 36461 15691
rect 36412 15660 36461 15688
rect 36412 15648 36418 15660
rect 36449 15657 36461 15660
rect 36495 15688 36507 15691
rect 36538 15688 36544 15700
rect 36495 15660 36544 15688
rect 36495 15657 36507 15660
rect 36449 15651 36507 15657
rect 36538 15648 36544 15660
rect 36596 15648 36602 15700
rect 41874 15648 41880 15700
rect 41932 15688 41938 15700
rect 41932 15660 44312 15688
rect 41932 15648 41938 15660
rect 21836 15592 24624 15620
rect 27709 15623 27767 15629
rect 13188 15524 15240 15552
rect 16945 15555 17003 15561
rect 9677 15487 9735 15493
rect 9677 15484 9689 15487
rect 9272 15456 9365 15484
rect 9416 15456 9689 15484
rect 9272 15444 9278 15456
rect 9677 15453 9689 15456
rect 9723 15453 9735 15487
rect 10410 15484 10416 15496
rect 10371 15456 10416 15484
rect 9677 15447 9735 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 12066 15484 12072 15496
rect 10928 15456 12072 15484
rect 10928 15444 10934 15456
rect 12066 15444 12072 15456
rect 12124 15484 12130 15496
rect 13188 15484 13216 15524
rect 16945 15521 16957 15555
rect 16991 15552 17003 15555
rect 18782 15552 18788 15564
rect 16991 15524 18788 15552
rect 16991 15521 17003 15524
rect 16945 15515 17003 15521
rect 18782 15512 18788 15524
rect 18840 15512 18846 15564
rect 20070 15552 20076 15564
rect 20031 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 21836 15561 21864 15592
rect 27709 15589 27721 15623
rect 27755 15620 27767 15623
rect 32030 15620 32036 15632
rect 27755 15592 32036 15620
rect 27755 15589 27767 15592
rect 27709 15583 27767 15589
rect 32030 15580 32036 15592
rect 32088 15580 32094 15632
rect 32125 15623 32183 15629
rect 32125 15589 32137 15623
rect 32171 15620 32183 15623
rect 32214 15620 32220 15632
rect 32171 15592 32220 15620
rect 32171 15589 32183 15592
rect 32125 15583 32183 15589
rect 32214 15580 32220 15592
rect 32272 15580 32278 15632
rect 33520 15592 34836 15620
rect 21821 15555 21879 15561
rect 21821 15521 21833 15555
rect 21867 15521 21879 15555
rect 24302 15552 24308 15564
rect 21821 15515 21879 15521
rect 22388 15524 24308 15552
rect 13354 15484 13360 15496
rect 12124 15456 13216 15484
rect 13315 15456 13360 15484
rect 12124 15444 12130 15456
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 15194 15484 15200 15496
rect 14507 15456 15200 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 15194 15444 15200 15456
rect 15252 15444 15258 15496
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15484 18107 15487
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 18095 15456 18521 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 18509 15453 18521 15456
rect 18555 15484 18567 15487
rect 19518 15484 19524 15496
rect 18555 15456 19524 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 19794 15484 19800 15496
rect 19755 15456 19800 15484
rect 19794 15444 19800 15456
rect 19852 15444 19858 15496
rect 22388 15493 22416 15524
rect 24302 15512 24308 15524
rect 24360 15512 24366 15564
rect 25409 15555 25467 15561
rect 25409 15521 25421 15555
rect 25455 15552 25467 15555
rect 25961 15555 26019 15561
rect 25961 15552 25973 15555
rect 25455 15524 25973 15552
rect 25455 15521 25467 15524
rect 25409 15515 25467 15521
rect 25961 15521 25973 15524
rect 26007 15521 26019 15555
rect 25961 15515 26019 15521
rect 26237 15555 26295 15561
rect 26237 15521 26249 15555
rect 26283 15552 26295 15555
rect 28905 15555 28963 15561
rect 28905 15552 28917 15555
rect 26283 15524 28917 15552
rect 26283 15521 26295 15524
rect 26237 15515 26295 15521
rect 28905 15521 28917 15524
rect 28951 15521 28963 15555
rect 29454 15552 29460 15564
rect 28905 15515 28963 15521
rect 29012 15524 29460 15552
rect 22373 15487 22431 15493
rect 21206 15456 22094 15484
rect 8662 15416 8668 15428
rect 5368 15388 8668 15416
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 11057 15419 11115 15425
rect 11057 15385 11069 15419
rect 11103 15385 11115 15419
rect 11057 15379 11115 15385
rect 5994 15348 6000 15360
rect 5955 15320 6000 15348
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 7558 15348 7564 15360
rect 7519 15320 7564 15348
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 10597 15351 10655 15357
rect 10597 15317 10609 15351
rect 10643 15348 10655 15351
rect 11072 15348 11100 15379
rect 13906 15376 13912 15428
rect 13964 15416 13970 15428
rect 16666 15416 16672 15428
rect 13964 15388 15502 15416
rect 16627 15388 16672 15416
rect 13964 15376 13970 15388
rect 16666 15376 16672 15388
rect 16724 15376 16730 15428
rect 22066 15416 22094 15456
rect 22373 15453 22385 15487
rect 22419 15453 22431 15487
rect 23014 15484 23020 15496
rect 22975 15456 23020 15484
rect 22373 15447 22431 15453
rect 23014 15444 23020 15456
rect 23072 15444 23078 15496
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15484 23719 15487
rect 24026 15484 24032 15496
rect 23707 15456 24032 15484
rect 23707 15453 23719 15456
rect 23661 15447 23719 15453
rect 24026 15444 24032 15456
rect 24084 15444 24090 15496
rect 24578 15484 24584 15496
rect 24539 15456 24584 15484
rect 24578 15444 24584 15456
rect 24636 15444 24642 15496
rect 25501 15487 25559 15493
rect 25501 15453 25513 15487
rect 25547 15453 25559 15487
rect 25501 15447 25559 15453
rect 22278 15416 22284 15428
rect 22066 15388 22284 15416
rect 22278 15376 22284 15388
rect 22336 15376 22342 15428
rect 22465 15419 22523 15425
rect 22465 15385 22477 15419
rect 22511 15416 22523 15419
rect 23474 15416 23480 15428
rect 22511 15388 23480 15416
rect 22511 15385 22523 15388
rect 22465 15379 22523 15385
rect 23474 15376 23480 15388
rect 23532 15376 23538 15428
rect 10643 15320 11100 15348
rect 13449 15351 13507 15357
rect 10643 15317 10655 15320
rect 10597 15311 10655 15317
rect 13449 15317 13461 15351
rect 13495 15348 13507 15351
rect 13814 15348 13820 15360
rect 13495 15320 13820 15348
rect 13495 15317 13507 15320
rect 13449 15311 13507 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 23201 15351 23259 15357
rect 23201 15317 23213 15351
rect 23247 15348 23259 15351
rect 24670 15348 24676 15360
rect 23247 15320 24676 15348
rect 23247 15317 23259 15320
rect 23201 15311 23259 15317
rect 24670 15308 24676 15320
rect 24728 15308 24734 15360
rect 25516 15348 25544 15447
rect 27522 15444 27528 15496
rect 27580 15484 27586 15496
rect 29012 15493 29040 15524
rect 29454 15512 29460 15524
rect 29512 15552 29518 15564
rect 33520 15552 33548 15592
rect 29512 15524 33548 15552
rect 29512 15512 29518 15524
rect 33594 15512 33600 15564
rect 33652 15552 33658 15564
rect 34701 15555 34759 15561
rect 34701 15552 34713 15555
rect 33652 15524 34713 15552
rect 33652 15512 33658 15524
rect 34701 15521 34713 15524
rect 34747 15521 34759 15555
rect 34808 15552 34836 15592
rect 36078 15580 36084 15632
rect 36136 15580 36142 15632
rect 39666 15620 39672 15632
rect 38764 15592 39672 15620
rect 36096 15552 36124 15580
rect 34808 15524 37136 15552
rect 34701 15515 34759 15521
rect 28169 15487 28227 15493
rect 28169 15484 28181 15487
rect 27580 15456 28181 15484
rect 27580 15444 27586 15456
rect 28169 15453 28181 15456
rect 28215 15453 28227 15487
rect 28169 15447 28227 15453
rect 28997 15487 29055 15493
rect 28997 15453 29009 15487
rect 29043 15453 29055 15487
rect 29546 15484 29552 15496
rect 29507 15456 29552 15484
rect 28997 15447 29055 15453
rect 29546 15444 29552 15456
rect 29604 15444 29610 15496
rect 33134 15484 33140 15496
rect 33095 15456 33140 15484
rect 33134 15444 33140 15456
rect 33192 15444 33198 15496
rect 33321 15487 33379 15493
rect 33321 15453 33333 15487
rect 33367 15484 33379 15487
rect 33873 15487 33931 15493
rect 33873 15484 33885 15487
rect 33367 15456 33885 15484
rect 33367 15453 33379 15456
rect 33321 15447 33379 15453
rect 33873 15453 33885 15456
rect 33919 15453 33931 15487
rect 33873 15447 33931 15453
rect 33962 15444 33968 15496
rect 34020 15484 34026 15496
rect 37108 15493 37136 15524
rect 38654 15512 38660 15564
rect 38712 15552 38718 15564
rect 38764 15561 38792 15592
rect 39666 15580 39672 15592
rect 39724 15580 39730 15632
rect 38749 15555 38807 15561
rect 38749 15552 38761 15555
rect 38712 15524 38761 15552
rect 38712 15512 38718 15524
rect 38749 15521 38761 15524
rect 38795 15521 38807 15555
rect 38749 15515 38807 15521
rect 38838 15512 38844 15564
rect 38896 15552 38902 15564
rect 39025 15555 39083 15561
rect 39025 15552 39037 15555
rect 38896 15524 39037 15552
rect 38896 15512 38902 15524
rect 39025 15521 39037 15524
rect 39071 15552 39083 15555
rect 39942 15552 39948 15564
rect 39071 15524 39948 15552
rect 39071 15521 39083 15524
rect 39025 15515 39083 15521
rect 39942 15512 39948 15524
rect 40000 15512 40006 15564
rect 40405 15555 40463 15561
rect 40405 15521 40417 15555
rect 40451 15552 40463 15555
rect 41601 15555 41659 15561
rect 41601 15552 41613 15555
rect 40451 15524 41613 15552
rect 40451 15521 40463 15524
rect 40405 15515 40463 15521
rect 41601 15521 41613 15524
rect 41647 15521 41659 15555
rect 41601 15515 41659 15521
rect 44177 15555 44235 15561
rect 44177 15521 44189 15555
rect 44223 15521 44235 15555
rect 44284 15552 44312 15660
rect 47670 15648 47676 15700
rect 47728 15688 47734 15700
rect 49694 15688 49700 15700
rect 47728 15660 49700 15688
rect 47728 15648 47734 15660
rect 49694 15648 49700 15660
rect 49752 15648 49758 15700
rect 51166 15688 51172 15700
rect 51127 15660 51172 15688
rect 51166 15648 51172 15660
rect 51224 15648 51230 15700
rect 53009 15691 53067 15697
rect 53009 15657 53021 15691
rect 53055 15688 53067 15691
rect 53374 15688 53380 15700
rect 53055 15660 53380 15688
rect 53055 15657 53067 15660
rect 53009 15651 53067 15657
rect 53374 15648 53380 15660
rect 53432 15648 53438 15700
rect 54113 15691 54171 15697
rect 54113 15657 54125 15691
rect 54159 15688 54171 15691
rect 54754 15688 54760 15700
rect 54159 15660 54760 15688
rect 54159 15657 54171 15660
rect 54113 15651 54171 15657
rect 54754 15648 54760 15660
rect 54812 15648 54818 15700
rect 55490 15648 55496 15700
rect 55548 15688 55554 15700
rect 58069 15691 58127 15697
rect 58069 15688 58081 15691
rect 55548 15660 58081 15688
rect 55548 15648 55554 15660
rect 58069 15657 58081 15660
rect 58115 15657 58127 15691
rect 58069 15651 58127 15657
rect 44453 15623 44511 15629
rect 44453 15589 44465 15623
rect 44499 15620 44511 15623
rect 44634 15620 44640 15632
rect 44499 15592 44640 15620
rect 44499 15589 44511 15592
rect 44453 15583 44511 15589
rect 44634 15580 44640 15592
rect 44692 15580 44698 15632
rect 48130 15580 48136 15632
rect 48188 15620 48194 15632
rect 54938 15620 54944 15632
rect 48188 15592 54944 15620
rect 48188 15580 48194 15592
rect 45189 15555 45247 15561
rect 45189 15552 45201 15555
rect 44284 15524 45201 15552
rect 44177 15515 44235 15521
rect 45189 15521 45201 15524
rect 45235 15521 45247 15555
rect 45922 15552 45928 15564
rect 45883 15524 45928 15552
rect 45189 15515 45247 15521
rect 37093 15487 37151 15493
rect 34020 15456 34065 15484
rect 34020 15444 34026 15456
rect 37093 15453 37105 15487
rect 37139 15453 37151 15487
rect 37642 15484 37648 15496
rect 37603 15456 37648 15484
rect 37093 15447 37151 15453
rect 37642 15444 37648 15456
rect 37700 15444 37706 15496
rect 38930 15444 38936 15496
rect 38988 15484 38994 15496
rect 39117 15487 39175 15493
rect 39117 15484 39129 15487
rect 38988 15456 39129 15484
rect 38988 15444 38994 15456
rect 39117 15453 39129 15456
rect 39163 15484 39175 15487
rect 40037 15487 40095 15493
rect 40037 15484 40049 15487
rect 39163 15456 40049 15484
rect 39163 15453 39175 15456
rect 39117 15447 39175 15453
rect 40037 15453 40049 15456
rect 40083 15453 40095 15487
rect 40862 15484 40868 15496
rect 40823 15456 40868 15484
rect 40037 15447 40095 15453
rect 40862 15444 40868 15456
rect 40920 15444 40926 15496
rect 44082 15484 44088 15496
rect 44043 15456 44088 15484
rect 44082 15444 44088 15456
rect 44140 15444 44146 15496
rect 27982 15416 27988 15428
rect 27462 15388 27988 15416
rect 27982 15376 27988 15388
rect 28040 15376 28046 15428
rect 29086 15376 29092 15428
rect 29144 15416 29150 15428
rect 29733 15419 29791 15425
rect 29733 15416 29745 15419
rect 29144 15388 29745 15416
rect 29144 15376 29150 15388
rect 29733 15385 29745 15388
rect 29779 15385 29791 15419
rect 31386 15416 31392 15428
rect 31347 15388 31392 15416
rect 29733 15379 29791 15385
rect 31386 15376 31392 15388
rect 31444 15416 31450 15428
rect 31570 15416 31576 15428
rect 31444 15388 31576 15416
rect 31444 15376 31450 15388
rect 31570 15376 31576 15388
rect 31628 15376 31634 15428
rect 32398 15376 32404 15428
rect 32456 15416 32462 15428
rect 34977 15419 35035 15425
rect 34977 15416 34989 15419
rect 32456 15388 34989 15416
rect 32456 15376 32462 15388
rect 34977 15385 34989 15388
rect 35023 15385 35035 15419
rect 34977 15379 35035 15385
rect 35250 15376 35256 15428
rect 35308 15416 35314 15428
rect 38378 15416 38384 15428
rect 35308 15388 35466 15416
rect 36372 15388 38384 15416
rect 35308 15376 35314 15388
rect 26602 15348 26608 15360
rect 25516 15320 26608 15348
rect 26602 15308 26608 15320
rect 26660 15308 26666 15360
rect 28810 15308 28816 15360
rect 28868 15348 28874 15360
rect 32214 15348 32220 15360
rect 28868 15320 32220 15348
rect 28868 15308 28874 15320
rect 32214 15308 32220 15320
rect 32272 15308 32278 15360
rect 33229 15351 33287 15357
rect 33229 15317 33241 15351
rect 33275 15348 33287 15351
rect 36372 15348 36400 15388
rect 38378 15376 38384 15388
rect 38436 15376 38442 15428
rect 41874 15416 41880 15428
rect 41835 15388 41880 15416
rect 41874 15376 41880 15388
rect 41932 15376 41938 15428
rect 44192 15416 44220 15515
rect 45922 15512 45928 15524
rect 45980 15512 45986 15564
rect 46014 15512 46020 15564
rect 46072 15552 46078 15564
rect 48222 15552 48228 15564
rect 46072 15524 46980 15552
rect 48183 15524 48228 15552
rect 46072 15512 46078 15524
rect 45002 15484 45008 15496
rect 44963 15456 45008 15484
rect 45002 15444 45008 15456
rect 45060 15444 45066 15496
rect 46952 15484 46980 15524
rect 48222 15512 48228 15524
rect 48280 15512 48286 15564
rect 49145 15555 49203 15561
rect 49145 15521 49157 15555
rect 49191 15552 49203 15555
rect 49234 15552 49240 15564
rect 49191 15524 49240 15552
rect 49191 15521 49203 15524
rect 49145 15515 49203 15521
rect 49234 15512 49240 15524
rect 49292 15512 49298 15564
rect 48395 15487 48453 15493
rect 46952 15456 48314 15484
rect 46106 15416 46112 15428
rect 41984 15388 42366 15416
rect 44192 15388 46112 15416
rect 33275 15320 36400 15348
rect 33275 15317 33287 15320
rect 33229 15311 33287 15317
rect 36538 15308 36544 15360
rect 36596 15348 36602 15360
rect 37001 15351 37059 15357
rect 37001 15348 37013 15351
rect 36596 15320 37013 15348
rect 36596 15308 36602 15320
rect 37001 15317 37013 15320
rect 37047 15317 37059 15351
rect 37001 15311 37059 15317
rect 37737 15351 37795 15357
rect 37737 15317 37749 15351
rect 37783 15348 37795 15351
rect 38746 15348 38752 15360
rect 37783 15320 38752 15348
rect 37783 15317 37795 15320
rect 37737 15311 37795 15317
rect 38746 15308 38752 15320
rect 38804 15308 38810 15360
rect 40957 15351 41015 15357
rect 40957 15317 40969 15351
rect 41003 15348 41015 15351
rect 41984 15348 42012 15388
rect 46106 15376 46112 15388
rect 46164 15376 46170 15428
rect 46934 15376 46940 15428
rect 46992 15416 46998 15428
rect 47486 15416 47492 15428
rect 46992 15388 47492 15416
rect 46992 15376 46998 15388
rect 47486 15376 47492 15388
rect 47544 15376 47550 15428
rect 48286 15416 48314 15456
rect 48395 15453 48407 15487
rect 48441 15484 48453 15487
rect 48441 15456 49372 15484
rect 48441 15453 48453 15456
rect 48395 15447 48453 15453
rect 49344 15428 49372 15456
rect 49786 15444 49792 15496
rect 49844 15484 49850 15496
rect 50157 15487 50215 15493
rect 50157 15484 50169 15487
rect 49844 15456 50169 15484
rect 49844 15444 49850 15456
rect 50157 15453 50169 15456
rect 50203 15453 50215 15487
rect 50157 15447 50215 15453
rect 51074 15444 51080 15496
rect 51132 15484 51138 15496
rect 51258 15484 51264 15496
rect 51132 15456 51177 15484
rect 51219 15456 51264 15484
rect 51132 15444 51138 15456
rect 51258 15444 51264 15456
rect 51316 15444 51322 15496
rect 51905 15487 51963 15493
rect 51905 15453 51917 15487
rect 51951 15484 51963 15487
rect 52104 15484 52132 15592
rect 54938 15580 54944 15592
rect 54996 15580 55002 15632
rect 52822 15512 52828 15564
rect 52880 15552 52886 15564
rect 54665 15555 54723 15561
rect 54665 15552 54677 15555
rect 52880 15524 54677 15552
rect 52880 15512 52886 15524
rect 54665 15521 54677 15524
rect 54711 15521 54723 15555
rect 56318 15552 56324 15564
rect 56279 15524 56324 15552
rect 54665 15515 54723 15521
rect 56318 15512 56324 15524
rect 56376 15512 56382 15564
rect 56594 15552 56600 15564
rect 56555 15524 56600 15552
rect 56594 15512 56600 15524
rect 56652 15512 56658 15564
rect 51951 15456 52132 15484
rect 51951 15453 51963 15456
rect 51905 15447 51963 15453
rect 52178 15444 52184 15496
rect 52236 15484 52242 15496
rect 53834 15484 53840 15496
rect 52236 15456 52281 15484
rect 52656 15456 53840 15484
rect 52236 15444 52242 15456
rect 49326 15416 49332 15428
rect 48286 15388 48820 15416
rect 49239 15388 49332 15416
rect 41003 15320 42012 15348
rect 43349 15351 43407 15357
rect 41003 15317 41015 15320
rect 40957 15311 41015 15317
rect 43349 15317 43361 15351
rect 43395 15348 43407 15351
rect 44634 15348 44640 15360
rect 43395 15320 44640 15348
rect 43395 15317 43407 15320
rect 43349 15311 43407 15317
rect 44634 15308 44640 15320
rect 44692 15308 44698 15360
rect 44818 15308 44824 15360
rect 44876 15348 44882 15360
rect 45922 15348 45928 15360
rect 44876 15320 45928 15348
rect 44876 15308 44882 15320
rect 45922 15308 45928 15320
rect 45980 15308 45986 15360
rect 47302 15308 47308 15360
rect 47360 15348 47366 15360
rect 47581 15351 47639 15357
rect 47581 15348 47593 15351
rect 47360 15320 47593 15348
rect 47360 15308 47366 15320
rect 47581 15317 47593 15320
rect 47627 15348 47639 15351
rect 48130 15348 48136 15360
rect 47627 15320 48136 15348
rect 47627 15317 47639 15320
rect 47581 15311 47639 15317
rect 48130 15308 48136 15320
rect 48188 15308 48194 15360
rect 48682 15348 48688 15360
rect 48643 15320 48688 15348
rect 48682 15308 48688 15320
rect 48740 15308 48746 15360
rect 48792 15348 48820 15388
rect 49326 15376 49332 15388
rect 49384 15416 49390 15428
rect 50706 15416 50712 15428
rect 49384 15388 50712 15416
rect 49384 15376 49390 15388
rect 50706 15376 50712 15388
rect 50764 15376 50770 15428
rect 52089 15419 52147 15425
rect 52089 15385 52101 15419
rect 52135 15416 52147 15419
rect 52656 15416 52684 15456
rect 53834 15444 53840 15456
rect 53892 15444 53898 15496
rect 53929 15487 53987 15493
rect 53929 15453 53941 15487
rect 53975 15453 53987 15487
rect 53929 15447 53987 15453
rect 54021 15487 54079 15493
rect 54021 15453 54033 15487
rect 54067 15484 54079 15487
rect 54110 15484 54116 15496
rect 54067 15456 54116 15484
rect 54067 15453 54079 15456
rect 54021 15447 54079 15453
rect 52135 15388 52684 15416
rect 52135 15385 52147 15388
rect 52089 15379 52147 15385
rect 52730 15376 52736 15428
rect 52788 15416 52794 15428
rect 52977 15419 53035 15425
rect 52977 15416 52989 15419
rect 52788 15388 52989 15416
rect 52788 15376 52794 15388
rect 52977 15385 52989 15388
rect 53023 15385 53035 15419
rect 53190 15416 53196 15428
rect 53151 15388 53196 15416
rect 52977 15379 53035 15385
rect 53190 15376 53196 15388
rect 53248 15376 53254 15428
rect 53558 15376 53564 15428
rect 53616 15416 53622 15428
rect 53944 15416 53972 15447
rect 54110 15444 54116 15456
rect 54168 15444 54174 15496
rect 54202 15444 54208 15496
rect 54260 15484 54266 15496
rect 55766 15484 55772 15496
rect 54260 15456 55772 15484
rect 54260 15444 54266 15456
rect 55766 15444 55772 15456
rect 55824 15444 55830 15496
rect 53616 15388 53972 15416
rect 53616 15376 53622 15388
rect 57330 15376 57336 15428
rect 57388 15376 57394 15428
rect 49234 15348 49240 15360
rect 48792 15320 49240 15348
rect 49234 15308 49240 15320
rect 49292 15308 49298 15360
rect 49970 15308 49976 15360
rect 50028 15348 50034 15360
rect 50341 15351 50399 15357
rect 50341 15348 50353 15351
rect 50028 15320 50353 15348
rect 50028 15308 50034 15320
rect 50341 15317 50353 15320
rect 50387 15317 50399 15351
rect 50341 15311 50399 15317
rect 51721 15351 51779 15357
rect 51721 15317 51733 15351
rect 51767 15348 51779 15351
rect 51902 15348 51908 15360
rect 51767 15320 51908 15348
rect 51767 15317 51779 15320
rect 51721 15311 51779 15317
rect 51902 15308 51908 15320
rect 51960 15308 51966 15360
rect 52822 15348 52828 15360
rect 52735 15320 52828 15348
rect 52822 15308 52828 15320
rect 52880 15348 52886 15360
rect 53650 15348 53656 15360
rect 52880 15320 53656 15348
rect 52880 15308 52886 15320
rect 53650 15308 53656 15320
rect 53708 15308 53714 15360
rect 1104 15258 58880 15280
rect 1104 15206 15398 15258
rect 15450 15206 15462 15258
rect 15514 15206 15526 15258
rect 15578 15206 15590 15258
rect 15642 15206 15654 15258
rect 15706 15206 29846 15258
rect 29898 15206 29910 15258
rect 29962 15206 29974 15258
rect 30026 15206 30038 15258
rect 30090 15206 30102 15258
rect 30154 15206 44294 15258
rect 44346 15206 44358 15258
rect 44410 15206 44422 15258
rect 44474 15206 44486 15258
rect 44538 15206 44550 15258
rect 44602 15206 58880 15258
rect 1104 15184 58880 15206
rect 5261 15147 5319 15153
rect 5261 15113 5273 15147
rect 5307 15144 5319 15147
rect 5350 15144 5356 15156
rect 5307 15116 5356 15144
rect 5307 15113 5319 15116
rect 5261 15107 5319 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 6822 15104 6828 15156
rect 6880 15144 6886 15156
rect 6880 15116 10732 15144
rect 6880 15104 6886 15116
rect 10704 15085 10732 15116
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 10928 15116 12434 15144
rect 10928 15104 10934 15116
rect 8665 15079 8723 15085
rect 8665 15045 8677 15079
rect 8711 15076 8723 15079
rect 10689 15079 10747 15085
rect 8711 15048 9522 15076
rect 8711 15045 8723 15048
rect 8665 15039 8723 15045
rect 10689 15045 10701 15079
rect 10735 15045 10747 15079
rect 12406 15076 12434 15116
rect 15194 15104 15200 15156
rect 15252 15144 15258 15156
rect 15657 15147 15715 15153
rect 15657 15144 15669 15147
rect 15252 15116 15669 15144
rect 15252 15104 15258 15116
rect 15657 15113 15669 15116
rect 15703 15113 15715 15147
rect 19426 15144 19432 15156
rect 15657 15107 15715 15113
rect 16592 15116 19432 15144
rect 12526 15076 12532 15088
rect 12406 15048 12532 15076
rect 10689 15039 10747 15045
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 14369 15079 14427 15085
rect 14369 15045 14381 15079
rect 14415 15076 14427 15079
rect 15286 15076 15292 15088
rect 14415 15048 15292 15076
rect 14415 15045 14427 15048
rect 14369 15039 14427 15045
rect 15286 15036 15292 15048
rect 15344 15036 15350 15088
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 5721 15011 5779 15017
rect 5721 15008 5733 15011
rect 5316 14980 5733 15008
rect 5316 14968 5322 14980
rect 5721 14977 5733 14980
rect 5767 14977 5779 15011
rect 5721 14971 5779 14977
rect 6362 14968 6368 15020
rect 6420 15008 6426 15020
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6420 14980 6653 15008
rect 6420 14968 6426 14980
rect 6641 14977 6653 14980
rect 6687 14977 6699 15011
rect 7466 15008 7472 15020
rect 7427 14980 7472 15008
rect 6641 14971 6699 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 7926 15008 7932 15020
rect 7887 14980 7932 15008
rect 7926 14968 7932 14980
rect 7984 15008 7990 15020
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 7984 14980 8585 15008
rect 7984 14968 7990 14980
rect 8573 14977 8585 14980
rect 8619 14977 8631 15011
rect 8573 14971 8631 14977
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 14977 11575 15011
rect 16592 15008 16620 15116
rect 19426 15104 19432 15116
rect 19484 15144 19490 15156
rect 20162 15144 20168 15156
rect 19484 15116 20168 15144
rect 19484 15104 19490 15116
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 21082 15144 21088 15156
rect 20640 15116 21088 15144
rect 16853 15079 16911 15085
rect 16853 15045 16865 15079
rect 16899 15076 16911 15079
rect 16899 15048 17802 15076
rect 16899 15045 16911 15048
rect 16853 15039 16911 15045
rect 19242 15036 19248 15088
rect 19300 15076 19306 15088
rect 20640 15076 20668 15116
rect 21082 15104 21088 15116
rect 21140 15104 21146 15156
rect 21269 15147 21327 15153
rect 21269 15113 21281 15147
rect 21315 15144 21327 15147
rect 21358 15144 21364 15156
rect 21315 15116 21364 15144
rect 21315 15113 21327 15116
rect 21269 15107 21327 15113
rect 21358 15104 21364 15116
rect 21416 15144 21422 15156
rect 21416 15116 26234 15144
rect 21416 15104 21422 15116
rect 19300 15048 20668 15076
rect 19300 15036 19306 15048
rect 20714 15036 20720 15088
rect 20772 15076 20778 15088
rect 21818 15076 21824 15088
rect 20772 15048 21824 15076
rect 20772 15036 20778 15048
rect 21818 15036 21824 15048
rect 21876 15036 21882 15088
rect 22186 15076 22192 15088
rect 22066 15048 22192 15076
rect 16758 15008 16764 15020
rect 13570 14980 16620 15008
rect 16719 14980 16764 15008
rect 11517 14971 11575 14977
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14940 7435 14943
rect 10594 14940 10600 14952
rect 7423 14912 10600 14940
rect 7423 14909 7435 14912
rect 7377 14903 7435 14909
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 10965 14943 11023 14949
rect 10965 14940 10977 14943
rect 10744 14912 10977 14940
rect 10744 14900 10750 14912
rect 10965 14909 10977 14912
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 6546 14832 6552 14884
rect 6604 14872 6610 14884
rect 9217 14875 9275 14881
rect 9217 14872 9229 14875
rect 6604 14844 9229 14872
rect 6604 14832 6610 14844
rect 9217 14841 9229 14844
rect 9263 14841 9275 14875
rect 9217 14835 9275 14841
rect 6733 14807 6791 14813
rect 6733 14773 6745 14807
rect 6779 14804 6791 14807
rect 7834 14804 7840 14816
rect 6779 14776 7840 14804
rect 6779 14773 6791 14776
rect 6733 14767 6791 14773
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 8018 14804 8024 14816
rect 7979 14776 8024 14804
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 11532 14804 11560 14971
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 15008 20683 15011
rect 20806 15008 20812 15020
rect 20671 14980 20812 15008
rect 20671 14977 20683 14980
rect 20625 14971 20683 14977
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 15008 20959 15011
rect 21082 15008 21088 15020
rect 20947 14980 21088 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 21082 14968 21088 14980
rect 21140 15008 21146 15020
rect 22066 15008 22094 15048
rect 22186 15036 22192 15048
rect 22244 15036 22250 15088
rect 24670 15076 24676 15088
rect 24631 15048 24676 15076
rect 24670 15036 24676 15048
rect 24728 15036 24734 15088
rect 26206 15076 26234 15116
rect 26970 15104 26976 15156
rect 27028 15144 27034 15156
rect 27433 15147 27491 15153
rect 27433 15144 27445 15147
rect 27028 15116 27445 15144
rect 27028 15104 27034 15116
rect 27433 15113 27445 15116
rect 27479 15144 27491 15147
rect 30466 15144 30472 15156
rect 27479 15116 30472 15144
rect 27479 15113 27491 15116
rect 27433 15107 27491 15113
rect 30466 15104 30472 15116
rect 30524 15144 30530 15156
rect 31205 15147 31263 15153
rect 31205 15144 31217 15147
rect 30524 15116 31217 15144
rect 30524 15104 30530 15116
rect 31205 15113 31217 15116
rect 31251 15113 31263 15147
rect 31205 15107 31263 15113
rect 32122 15104 32128 15156
rect 32180 15144 32186 15156
rect 32769 15147 32827 15153
rect 32769 15144 32781 15147
rect 32180 15116 32781 15144
rect 32180 15104 32186 15116
rect 32769 15113 32781 15116
rect 32815 15113 32827 15147
rect 32769 15107 32827 15113
rect 35158 15104 35164 15156
rect 35216 15144 35222 15156
rect 35345 15147 35403 15153
rect 35345 15144 35357 15147
rect 35216 15116 35357 15144
rect 35216 15104 35222 15116
rect 35345 15113 35357 15116
rect 35391 15144 35403 15147
rect 35434 15144 35440 15156
rect 35391 15116 35440 15144
rect 35391 15113 35403 15116
rect 35345 15107 35403 15113
rect 35434 15104 35440 15116
rect 35492 15104 35498 15156
rect 35986 15144 35992 15156
rect 35947 15116 35992 15144
rect 35986 15104 35992 15116
rect 36044 15104 36050 15156
rect 39577 15147 39635 15153
rect 39577 15144 39589 15147
rect 38580 15116 39589 15144
rect 27798 15076 27804 15088
rect 26206 15048 27804 15076
rect 24026 15008 24032 15020
rect 21140 14980 22094 15008
rect 23987 14980 24032 15008
rect 21140 14968 21146 14980
rect 24026 14968 24032 14980
rect 24084 14968 24090 15020
rect 27356 15017 27384 15048
rect 27798 15036 27804 15048
rect 27856 15076 27862 15088
rect 28626 15076 28632 15088
rect 27856 15048 28632 15076
rect 27856 15036 27862 15048
rect 28626 15036 28632 15048
rect 28684 15036 28690 15088
rect 30558 15076 30564 15088
rect 30519 15048 30564 15076
rect 30558 15036 30564 15048
rect 30616 15036 30622 15088
rect 35250 15076 35256 15088
rect 35098 15048 35256 15076
rect 35250 15036 35256 15048
rect 35308 15036 35314 15088
rect 38580 15076 38608 15116
rect 39577 15113 39589 15116
rect 39623 15113 39635 15147
rect 39577 15107 39635 15113
rect 39942 15104 39948 15156
rect 40000 15144 40006 15156
rect 40129 15147 40187 15153
rect 40129 15144 40141 15147
rect 40000 15116 40141 15144
rect 40000 15104 40006 15116
rect 40129 15113 40141 15116
rect 40175 15113 40187 15147
rect 40678 15144 40684 15156
rect 40129 15107 40187 15113
rect 40236 15116 40684 15144
rect 38746 15076 38752 15088
rect 38318 15048 38608 15076
rect 38707 15048 38752 15076
rect 38746 15036 38752 15048
rect 38804 15036 38810 15088
rect 27341 15011 27399 15017
rect 27341 14977 27353 15011
rect 27387 14977 27399 15011
rect 27341 14971 27399 14977
rect 27614 14968 27620 15020
rect 27672 15008 27678 15020
rect 27985 15011 28043 15017
rect 27985 15008 27997 15011
rect 27672 14980 27997 15008
rect 27672 14968 27678 14980
rect 27985 14977 27997 14980
rect 28031 14977 28043 15011
rect 32306 15008 32312 15020
rect 32267 14980 32312 15008
rect 27985 14971 28043 14977
rect 32306 14968 32312 14980
rect 32364 14968 32370 15020
rect 33594 15008 33600 15020
rect 33555 14980 33600 15008
rect 33594 14968 33600 14980
rect 33652 14968 33658 15020
rect 36081 15011 36139 15017
rect 36081 14977 36093 15011
rect 36127 15008 36139 15011
rect 36446 15008 36452 15020
rect 36127 14980 36452 15008
rect 36127 14977 36139 14980
rect 36081 14971 36139 14977
rect 36446 14968 36452 14980
rect 36504 14968 36510 15020
rect 36725 15011 36783 15017
rect 36725 14977 36737 15011
rect 36771 15008 36783 15011
rect 36771 14980 37320 15008
rect 36771 14977 36783 14980
rect 36725 14971 36783 14977
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 11655 14912 12173 14940
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 12161 14909 12173 14912
rect 12207 14909 12219 14943
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12161 14903 12219 14909
rect 12268 14912 12449 14940
rect 12268 14816 12296 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12526 14900 12532 14952
rect 12584 14940 12590 14952
rect 17494 14940 17500 14952
rect 12584 14912 14136 14940
rect 17455 14912 17500 14940
rect 12584 14900 12590 14912
rect 9732 14776 11560 14804
rect 9732 14764 9738 14776
rect 12250 14764 12256 14816
rect 12308 14764 12314 14816
rect 13909 14807 13967 14813
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 13998 14804 14004 14816
rect 13955 14776 14004 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14108 14804 14136 14912
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 18966 14940 18972 14952
rect 18927 14912 18972 14940
rect 18966 14900 18972 14912
rect 19024 14900 19030 14952
rect 19245 14943 19303 14949
rect 19245 14909 19257 14943
rect 19291 14940 19303 14943
rect 19702 14940 19708 14952
rect 19291 14912 19708 14940
rect 19291 14909 19303 14912
rect 19245 14903 19303 14909
rect 19702 14900 19708 14912
rect 19760 14940 19766 14952
rect 21634 14940 21640 14952
rect 19760 14912 21640 14940
rect 19760 14900 19766 14912
rect 21634 14900 21640 14912
rect 21692 14900 21698 14952
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 21968 14912 23244 14940
rect 21968 14900 21974 14912
rect 19518 14832 19524 14884
rect 19576 14872 19582 14884
rect 23109 14875 23167 14881
rect 23109 14872 23121 14875
rect 19576 14844 23121 14872
rect 19576 14832 19582 14844
rect 23109 14841 23121 14844
rect 23155 14841 23167 14875
rect 23216 14872 23244 14912
rect 23566 14900 23572 14952
rect 23624 14940 23630 14952
rect 28997 14943 29055 14949
rect 28997 14940 29009 14943
rect 23624 14912 29009 14940
rect 23624 14900 23630 14912
rect 28997 14909 29009 14912
rect 29043 14940 29055 14943
rect 29086 14940 29092 14952
rect 29043 14912 29092 14940
rect 29043 14909 29055 14912
rect 28997 14903 29055 14909
rect 29086 14900 29092 14912
rect 29144 14900 29150 14952
rect 30745 14943 30803 14949
rect 30745 14909 30757 14943
rect 30791 14940 30803 14943
rect 33042 14940 33048 14952
rect 30791 14912 33048 14940
rect 30791 14909 30803 14912
rect 30745 14903 30803 14909
rect 33042 14900 33048 14912
rect 33100 14900 33106 14952
rect 33226 14900 33232 14952
rect 33284 14940 33290 14952
rect 33873 14943 33931 14949
rect 33873 14940 33885 14943
rect 33284 14912 33885 14940
rect 33284 14900 33290 14912
rect 33873 14909 33885 14912
rect 33919 14909 33931 14943
rect 33873 14903 33931 14909
rect 26970 14872 26976 14884
rect 23216 14844 26976 14872
rect 23109 14835 23167 14841
rect 26970 14832 26976 14844
rect 27028 14832 27034 14884
rect 19886 14804 19892 14816
rect 14108 14776 19892 14804
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 24210 14804 24216 14816
rect 24171 14776 24216 14804
rect 24210 14764 24216 14776
rect 24268 14764 24274 14816
rect 25958 14804 25964 14816
rect 25919 14776 25964 14804
rect 25958 14764 25964 14776
rect 26016 14764 26022 14816
rect 28074 14804 28080 14816
rect 28035 14776 28080 14804
rect 28074 14764 28080 14776
rect 28132 14764 28138 14816
rect 32214 14804 32220 14816
rect 32175 14776 32220 14804
rect 32214 14764 32220 14776
rect 32272 14764 32278 14816
rect 36630 14804 36636 14816
rect 36591 14776 36636 14804
rect 36630 14764 36636 14776
rect 36688 14764 36694 14816
rect 37292 14813 37320 14980
rect 39022 14968 39028 15020
rect 39080 15008 39086 15020
rect 39669 15011 39727 15017
rect 39080 14980 39125 15008
rect 39080 14968 39086 14980
rect 39669 14977 39681 15011
rect 39715 15008 39727 15011
rect 40126 15008 40132 15020
rect 39715 14980 40132 15008
rect 39715 14977 39727 14980
rect 39669 14971 39727 14977
rect 40126 14968 40132 14980
rect 40184 15008 40190 15020
rect 40236 15008 40264 15116
rect 40678 15104 40684 15116
rect 40736 15104 40742 15156
rect 45002 15104 45008 15156
rect 45060 15144 45066 15156
rect 45462 15144 45468 15156
rect 45060 15116 45468 15144
rect 45060 15104 45066 15116
rect 45462 15104 45468 15116
rect 45520 15144 45526 15156
rect 50706 15144 50712 15156
rect 45520 15116 47900 15144
rect 50667 15116 50712 15144
rect 45520 15104 45526 15116
rect 41414 15076 41420 15088
rect 40184 14980 40264 15008
rect 40696 15048 41420 15076
rect 40184 14968 40190 14980
rect 40494 14900 40500 14952
rect 40552 14940 40558 14952
rect 40696 14949 40724 15048
rect 41414 15036 41420 15048
rect 41472 15036 41478 15088
rect 41874 15036 41880 15088
rect 41932 15076 41938 15088
rect 42429 15079 42487 15085
rect 42429 15076 42441 15079
rect 41932 15048 42441 15076
rect 41932 15036 41938 15048
rect 42429 15045 42441 15048
rect 42475 15045 42487 15079
rect 44726 15076 44732 15088
rect 42429 15039 42487 15045
rect 42720 15048 44732 15076
rect 40957 15011 41015 15017
rect 40957 14977 40969 15011
rect 41003 15008 41015 15011
rect 41138 15008 41144 15020
rect 41003 14980 41144 15008
rect 41003 14977 41015 14980
rect 40957 14971 41015 14977
rect 41138 14968 41144 14980
rect 41196 14968 41202 15020
rect 41693 15011 41751 15017
rect 41693 14977 41705 15011
rect 41739 15008 41751 15011
rect 41782 15008 41788 15020
rect 41739 14980 41788 15008
rect 41739 14977 41751 14980
rect 41693 14971 41751 14977
rect 41782 14968 41788 14980
rect 41840 14968 41846 15020
rect 42720 15017 42748 15048
rect 44726 15036 44732 15048
rect 44784 15076 44790 15088
rect 44784 15048 46060 15076
rect 44784 15036 44790 15048
rect 46032 15017 46060 15048
rect 46842 15036 46848 15088
rect 46900 15076 46906 15088
rect 46900 15048 47808 15076
rect 46900 15036 46906 15048
rect 42705 15011 42763 15017
rect 42705 14977 42717 15011
rect 42751 14977 42763 15011
rect 42705 14971 42763 14977
rect 46017 15011 46075 15017
rect 46017 14977 46029 15011
rect 46063 14977 46075 15011
rect 46017 14971 46075 14977
rect 47486 14968 47492 15020
rect 47544 15008 47550 15020
rect 47581 15011 47639 15017
rect 47581 15008 47593 15011
rect 47544 14980 47593 15008
rect 47544 14968 47550 14980
rect 47581 14977 47593 14980
rect 47627 14977 47639 15011
rect 47581 14971 47639 14977
rect 40681 14943 40739 14949
rect 40681 14940 40693 14943
rect 40552 14912 40693 14940
rect 40552 14900 40558 14912
rect 40681 14909 40693 14912
rect 40727 14909 40739 14943
rect 40681 14903 40739 14909
rect 41414 14900 41420 14952
rect 41472 14940 41478 14952
rect 42610 14940 42616 14952
rect 41472 14912 42616 14940
rect 41472 14900 41478 14912
rect 42610 14900 42616 14912
rect 42668 14940 42674 14952
rect 42886 14940 42892 14952
rect 42668 14912 42892 14940
rect 42668 14900 42674 14912
rect 42886 14900 42892 14912
rect 42944 14940 42950 14952
rect 44818 14940 44824 14952
rect 42944 14912 44824 14940
rect 42944 14900 42950 14912
rect 44818 14900 44824 14912
rect 44876 14900 44882 14952
rect 45094 14940 45100 14952
rect 45055 14912 45100 14940
rect 45094 14900 45100 14912
rect 45152 14900 45158 14952
rect 45281 14943 45339 14949
rect 45281 14909 45293 14943
rect 45327 14940 45339 14943
rect 45830 14940 45836 14952
rect 45327 14912 45836 14940
rect 45327 14909 45339 14912
rect 45281 14903 45339 14909
rect 45830 14900 45836 14912
rect 45888 14900 45894 14952
rect 47780 14949 47808 15048
rect 47872 15017 47900 15116
rect 50706 15104 50712 15116
rect 50764 15104 50770 15156
rect 52178 15104 52184 15156
rect 52236 15144 52242 15156
rect 52733 15147 52791 15153
rect 52733 15144 52745 15147
rect 52236 15116 52745 15144
rect 52236 15104 52242 15116
rect 52733 15113 52745 15116
rect 52779 15113 52791 15147
rect 55125 15147 55183 15153
rect 55125 15144 55137 15147
rect 52733 15107 52791 15113
rect 54312 15116 55137 15144
rect 48682 15036 48688 15088
rect 48740 15076 48746 15088
rect 49237 15079 49295 15085
rect 49237 15076 49249 15079
rect 48740 15048 49249 15076
rect 48740 15036 48746 15048
rect 49237 15045 49249 15048
rect 49283 15045 49295 15079
rect 49237 15039 49295 15045
rect 50246 15036 50252 15088
rect 50304 15036 50310 15088
rect 52822 15076 52828 15088
rect 51368 15048 52828 15076
rect 51368 15020 51396 15048
rect 52822 15036 52828 15048
rect 52880 15036 52886 15088
rect 54312 15076 54340 15116
rect 55125 15113 55137 15116
rect 55171 15113 55183 15147
rect 55125 15107 55183 15113
rect 53116 15048 54340 15076
rect 53116 15020 53144 15048
rect 47857 15011 47915 15017
rect 47857 14977 47869 15011
rect 47903 14977 47915 15011
rect 51350 15008 51356 15020
rect 51263 14980 51356 15008
rect 47857 14971 47915 14977
rect 51350 14968 51356 14980
rect 51408 14968 51414 15020
rect 51537 15011 51595 15017
rect 51537 14977 51549 15011
rect 51583 15008 51595 15011
rect 52917 15011 52975 15017
rect 51583 14980 51764 15008
rect 51583 14977 51595 14980
rect 51537 14971 51595 14977
rect 45925 14943 45983 14949
rect 45925 14909 45937 14943
rect 45971 14909 45983 14943
rect 45925 14903 45983 14909
rect 46845 14943 46903 14949
rect 46845 14909 46857 14943
rect 46891 14909 46903 14943
rect 46845 14903 46903 14909
rect 47765 14943 47823 14949
rect 47765 14909 47777 14943
rect 47811 14940 47823 14943
rect 48222 14940 48228 14952
rect 47811 14912 48228 14940
rect 47811 14909 47823 14912
rect 47765 14903 47823 14909
rect 44634 14832 44640 14884
rect 44692 14872 44698 14884
rect 45940 14872 45968 14903
rect 46860 14872 46888 14903
rect 48222 14900 48228 14912
rect 48280 14900 48286 14952
rect 48961 14943 49019 14949
rect 48961 14909 48973 14943
rect 49007 14940 49019 14943
rect 49786 14940 49792 14952
rect 49007 14912 49792 14940
rect 49007 14909 49019 14912
rect 48961 14903 49019 14909
rect 49786 14900 49792 14912
rect 49844 14900 49850 14952
rect 51442 14900 51448 14952
rect 51500 14940 51506 14952
rect 51629 14943 51687 14949
rect 51500 14912 51545 14940
rect 51500 14900 51506 14912
rect 51629 14909 51641 14943
rect 51675 14909 51687 14943
rect 51736 14940 51764 14980
rect 52917 14977 52929 15011
rect 52963 15008 52975 15011
rect 53098 15008 53104 15020
rect 52963 14980 53104 15008
rect 52963 14977 52975 14980
rect 52917 14971 52975 14977
rect 53098 14968 53104 14980
rect 53156 14968 53162 15020
rect 53193 15011 53251 15017
rect 53193 14977 53205 15011
rect 53239 15008 53251 15011
rect 53282 15008 53288 15020
rect 53239 14980 53288 15008
rect 53239 14977 53251 14980
rect 53193 14971 53251 14977
rect 53282 14968 53288 14980
rect 53340 14968 53346 15020
rect 54312 15017 54340 15048
rect 56042 15036 56048 15088
rect 56100 15036 56106 15088
rect 54297 15011 54355 15017
rect 54297 14977 54309 15011
rect 54343 14977 54355 15011
rect 54297 14971 54355 14977
rect 53009 14943 53067 14949
rect 53009 14940 53021 14943
rect 51736 14912 53021 14940
rect 51629 14903 51687 14909
rect 53009 14909 53021 14912
rect 53055 14940 53067 14943
rect 53466 14940 53472 14952
rect 53055 14912 53472 14940
rect 53055 14909 53067 14912
rect 53009 14903 53067 14909
rect 48866 14872 48872 14884
rect 44692 14844 45968 14872
rect 46124 14844 46520 14872
rect 46860 14844 48872 14872
rect 44692 14832 44698 14844
rect 37277 14807 37335 14813
rect 37277 14773 37289 14807
rect 37323 14804 37335 14807
rect 38286 14804 38292 14816
rect 37323 14776 38292 14804
rect 37323 14773 37335 14776
rect 37277 14767 37335 14773
rect 38286 14764 38292 14776
rect 38344 14764 38350 14816
rect 41877 14807 41935 14813
rect 41877 14773 41889 14807
rect 41923 14804 41935 14807
rect 42978 14804 42984 14816
rect 41923 14776 42984 14804
rect 41923 14773 41935 14776
rect 41877 14767 41935 14773
rect 42978 14764 42984 14776
rect 43036 14764 43042 14816
rect 44910 14764 44916 14816
rect 44968 14804 44974 14816
rect 46124 14804 46152 14844
rect 44968 14776 46152 14804
rect 46492 14804 46520 14844
rect 48866 14832 48872 14844
rect 48924 14832 48930 14884
rect 47581 14807 47639 14813
rect 47581 14804 47593 14807
rect 46492 14776 47593 14804
rect 44968 14764 44974 14776
rect 47581 14773 47593 14776
rect 47627 14773 47639 14807
rect 48038 14804 48044 14816
rect 47999 14776 48044 14804
rect 47581 14767 47639 14773
rect 48038 14764 48044 14776
rect 48096 14764 48102 14816
rect 49694 14764 49700 14816
rect 49752 14804 49758 14816
rect 51169 14807 51227 14813
rect 51169 14804 51181 14807
rect 49752 14776 51181 14804
rect 49752 14764 49758 14776
rect 51169 14773 51181 14776
rect 51215 14773 51227 14807
rect 51169 14767 51227 14773
rect 51258 14764 51264 14816
rect 51316 14804 51322 14816
rect 51644 14804 51672 14903
rect 53466 14900 53472 14912
rect 53524 14900 53530 14952
rect 53742 14900 53748 14952
rect 53800 14940 53806 14952
rect 54205 14943 54263 14949
rect 54205 14940 54217 14943
rect 53800 14912 54217 14940
rect 53800 14900 53806 14912
rect 54205 14909 54217 14912
rect 54251 14909 54263 14943
rect 56597 14943 56655 14949
rect 56597 14940 56609 14943
rect 54205 14903 54263 14909
rect 54680 14912 56609 14940
rect 54680 14881 54708 14912
rect 56597 14909 56609 14912
rect 56643 14909 56655 14943
rect 56870 14940 56876 14952
rect 56831 14912 56876 14940
rect 56597 14903 56655 14909
rect 56870 14900 56876 14912
rect 56928 14900 56934 14952
rect 54665 14875 54723 14881
rect 54665 14841 54677 14875
rect 54711 14841 54723 14875
rect 54665 14835 54723 14841
rect 51316 14776 51672 14804
rect 53193 14807 53251 14813
rect 51316 14764 51322 14776
rect 53193 14773 53205 14807
rect 53239 14804 53251 14807
rect 53374 14804 53380 14816
rect 53239 14776 53380 14804
rect 53239 14773 53251 14776
rect 53193 14767 53251 14773
rect 53374 14764 53380 14776
rect 53432 14804 53438 14816
rect 57146 14804 57152 14816
rect 53432 14776 57152 14804
rect 53432 14764 53438 14776
rect 57146 14764 57152 14776
rect 57204 14764 57210 14816
rect 1104 14714 58880 14736
rect 1104 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 8302 14714
rect 8354 14662 8366 14714
rect 8418 14662 8430 14714
rect 8482 14662 22622 14714
rect 22674 14662 22686 14714
rect 22738 14662 22750 14714
rect 22802 14662 22814 14714
rect 22866 14662 22878 14714
rect 22930 14662 37070 14714
rect 37122 14662 37134 14714
rect 37186 14662 37198 14714
rect 37250 14662 37262 14714
rect 37314 14662 37326 14714
rect 37378 14662 51518 14714
rect 51570 14662 51582 14714
rect 51634 14662 51646 14714
rect 51698 14662 51710 14714
rect 51762 14662 51774 14714
rect 51826 14662 58880 14714
rect 1104 14640 58880 14662
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5905 14603 5963 14609
rect 5905 14600 5917 14603
rect 5316 14572 5917 14600
rect 5316 14560 5322 14572
rect 5905 14569 5917 14572
rect 5951 14569 5963 14603
rect 5905 14563 5963 14569
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 6638 14600 6644 14612
rect 6595 14572 6644 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 7653 14603 7711 14609
rect 7653 14569 7665 14603
rect 7699 14600 7711 14603
rect 8846 14600 8852 14612
rect 7699 14572 8852 14600
rect 7699 14569 7711 14572
rect 7653 14563 7711 14569
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9861 14603 9919 14609
rect 9861 14569 9873 14603
rect 9907 14600 9919 14603
rect 9950 14600 9956 14612
rect 9907 14572 9956 14600
rect 9907 14569 9919 14572
rect 9861 14563 9919 14569
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10594 14560 10600 14612
rect 10652 14600 10658 14612
rect 11897 14603 11955 14609
rect 11897 14600 11909 14603
rect 10652 14572 11909 14600
rect 10652 14560 10658 14572
rect 11897 14569 11909 14572
rect 11943 14569 11955 14603
rect 11897 14563 11955 14569
rect 13449 14603 13507 14609
rect 13449 14569 13461 14603
rect 13495 14600 13507 14603
rect 13906 14600 13912 14612
rect 13495 14572 13912 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14734 14560 14740 14612
rect 14792 14600 14798 14612
rect 19242 14600 19248 14612
rect 14792 14572 19248 14600
rect 14792 14560 14798 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19613 14603 19671 14609
rect 19613 14569 19625 14603
rect 19659 14600 19671 14603
rect 19794 14600 19800 14612
rect 19659 14572 19800 14600
rect 19659 14569 19671 14572
rect 19613 14563 19671 14569
rect 19794 14560 19800 14572
rect 19852 14560 19858 14612
rect 19886 14560 19892 14612
rect 19944 14600 19950 14612
rect 23566 14600 23572 14612
rect 19944 14572 23572 14600
rect 19944 14560 19950 14572
rect 23566 14560 23572 14572
rect 23624 14560 23630 14612
rect 24762 14600 24768 14612
rect 24412 14572 24768 14600
rect 8294 14532 8300 14544
rect 8255 14504 8300 14532
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 8938 14492 8944 14544
rect 8996 14532 9002 14544
rect 10870 14532 10876 14544
rect 8996 14504 10876 14532
rect 8996 14492 9002 14504
rect 10870 14492 10876 14504
rect 10928 14492 10934 14544
rect 12897 14535 12955 14541
rect 12897 14501 12909 14535
rect 12943 14532 12955 14535
rect 14366 14532 14372 14544
rect 12943 14504 14372 14532
rect 12943 14501 12955 14504
rect 12897 14495 12955 14501
rect 14366 14492 14372 14504
rect 14424 14492 14430 14544
rect 19334 14492 19340 14544
rect 19392 14532 19398 14544
rect 20349 14535 20407 14541
rect 20349 14532 20361 14535
rect 19392 14504 20361 14532
rect 19392 14492 19398 14504
rect 20349 14501 20361 14504
rect 20395 14501 20407 14535
rect 20349 14495 20407 14501
rect 20456 14504 22232 14532
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 5960 14436 7604 14464
rect 5960 14424 5966 14436
rect 7576 14405 7604 14436
rect 7926 14424 7932 14476
rect 7984 14464 7990 14476
rect 7984 14436 9812 14464
rect 7984 14424 7990 14436
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14396 8263 14399
rect 8662 14396 8668 14408
rect 8251 14368 8668 14396
rect 8251 14365 8263 14368
rect 8205 14359 8263 14365
rect 6656 14328 6684 14359
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 9309 14399 9367 14405
rect 9309 14365 9321 14399
rect 9355 14396 9367 14399
rect 9674 14396 9680 14408
rect 9355 14368 9680 14396
rect 9355 14365 9367 14368
rect 9309 14359 9367 14365
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 9784 14405 9812 14436
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 14277 14467 14335 14473
rect 9916 14436 12756 14464
rect 9916 14424 9922 14436
rect 12728 14405 12756 14436
rect 14277 14433 14289 14467
rect 14323 14464 14335 14467
rect 15746 14464 15752 14476
rect 14323 14436 15752 14464
rect 14323 14433 14335 14436
rect 14277 14427 14335 14433
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 18506 14464 18512 14476
rect 16132 14436 18512 14464
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14365 9827 14399
rect 9769 14359 9827 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14396 12771 14399
rect 12802 14396 12808 14408
rect 12759 14368 12808 14396
rect 12759 14365 12771 14368
rect 12713 14359 12771 14365
rect 9217 14331 9275 14337
rect 6656 14300 7788 14328
rect 7760 14272 7788 14300
rect 9217 14297 9229 14331
rect 9263 14328 9275 14331
rect 9263 14300 10718 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 10413 14263 10471 14269
rect 10413 14260 10425 14263
rect 7800 14232 10425 14260
rect 7800 14220 7806 14232
rect 10413 14229 10425 14232
rect 10459 14229 10471 14263
rect 10413 14223 10471 14229
rect 10594 14220 10600 14272
rect 10652 14260 10658 14272
rect 12176 14260 12204 14359
rect 12802 14356 12808 14368
rect 12860 14356 12866 14408
rect 13354 14396 13360 14408
rect 13315 14368 13360 14396
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 16022 14356 16028 14408
rect 16080 14396 16086 14408
rect 16132 14396 16160 14436
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 16482 14396 16488 14408
rect 16080 14368 16173 14396
rect 16443 14368 16488 14396
rect 16080 14356 16086 14368
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 17126 14356 17132 14408
rect 17184 14396 17190 14408
rect 19518 14396 19524 14408
rect 17184 14368 19380 14396
rect 19479 14368 19524 14396
rect 17184 14356 17190 14368
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 13372 14328 13400 14356
rect 12492 14300 13400 14328
rect 12492 14288 12498 14300
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 15749 14331 15807 14337
rect 13872 14300 14582 14328
rect 13872 14288 13878 14300
rect 15749 14297 15761 14331
rect 15795 14328 15807 14331
rect 17310 14328 17316 14340
rect 15795 14300 17316 14328
rect 15795 14297 15807 14300
rect 15749 14291 15807 14297
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 19352 14328 19380 14368
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 20456 14405 20484 14504
rect 21174 14464 21180 14476
rect 21135 14436 21180 14464
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 22204 14464 22232 14504
rect 23934 14464 23940 14476
rect 22204 14436 23940 14464
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 24412 14473 24440 14572
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 27338 14560 27344 14612
rect 27396 14600 27402 14612
rect 28994 14600 29000 14612
rect 27396 14572 27752 14600
rect 28955 14572 29000 14600
rect 27396 14560 27402 14572
rect 26145 14535 26203 14541
rect 26145 14501 26157 14535
rect 26191 14532 26203 14535
rect 27614 14532 27620 14544
rect 26191 14504 27620 14532
rect 26191 14501 26203 14504
rect 26145 14495 26203 14501
rect 27614 14492 27620 14504
rect 27672 14492 27678 14544
rect 27724 14532 27752 14572
rect 28994 14560 29000 14572
rect 29052 14560 29058 14612
rect 33873 14603 33931 14609
rect 33873 14569 33885 14603
rect 33919 14600 33931 14603
rect 33962 14600 33968 14612
rect 33919 14572 33968 14600
rect 33919 14569 33931 14572
rect 33873 14563 33931 14569
rect 33962 14560 33968 14572
rect 34020 14560 34026 14612
rect 37090 14600 37096 14612
rect 35636 14572 37096 14600
rect 32306 14532 32312 14544
rect 27724 14504 30696 14532
rect 24397 14467 24455 14473
rect 24397 14433 24409 14467
rect 24443 14433 24455 14467
rect 24397 14427 24455 14433
rect 24673 14467 24731 14473
rect 24673 14433 24685 14467
rect 24719 14464 24731 14467
rect 28074 14464 28080 14476
rect 24719 14436 28080 14464
rect 24719 14433 24731 14436
rect 24673 14427 24731 14433
rect 28074 14424 28080 14436
rect 28132 14424 28138 14476
rect 30466 14424 30472 14476
rect 30524 14464 30530 14476
rect 30561 14467 30619 14473
rect 30561 14464 30573 14467
rect 30524 14436 30573 14464
rect 30524 14424 30530 14436
rect 30561 14433 30573 14436
rect 30607 14433 30619 14467
rect 30668 14464 30696 14504
rect 31864 14504 32312 14532
rect 31864 14464 31892 14504
rect 32306 14492 32312 14504
rect 32364 14532 32370 14544
rect 32861 14535 32919 14541
rect 32861 14532 32873 14535
rect 32364 14504 32873 14532
rect 32364 14492 32370 14504
rect 32861 14501 32873 14504
rect 32907 14532 32919 14535
rect 35636 14532 35664 14572
rect 37090 14560 37096 14572
rect 37148 14560 37154 14612
rect 45094 14600 45100 14612
rect 39132 14572 45100 14600
rect 32907 14504 35664 14532
rect 32907 14501 32919 14504
rect 32861 14495 32919 14501
rect 36630 14464 36636 14476
rect 30668 14436 31892 14464
rect 36591 14436 36636 14464
rect 30561 14427 30619 14433
rect 36630 14424 36636 14436
rect 36688 14424 36694 14476
rect 36909 14467 36967 14473
rect 36909 14433 36921 14467
rect 36955 14464 36967 14467
rect 38654 14464 38660 14476
rect 36955 14436 38660 14464
rect 36955 14433 36967 14436
rect 36909 14427 36967 14433
rect 38654 14424 38660 14436
rect 38712 14424 38718 14476
rect 39132 14473 39160 14572
rect 45094 14560 45100 14572
rect 45152 14560 45158 14612
rect 46106 14600 46112 14612
rect 46067 14572 46112 14600
rect 46106 14560 46112 14572
rect 46164 14560 46170 14612
rect 48501 14603 48559 14609
rect 48501 14569 48513 14603
rect 48547 14600 48559 14603
rect 48774 14600 48780 14612
rect 48547 14572 48780 14600
rect 48547 14569 48559 14572
rect 48501 14563 48559 14569
rect 48774 14560 48780 14572
rect 48832 14560 48838 14612
rect 48866 14560 48872 14612
rect 48924 14600 48930 14612
rect 52914 14600 52920 14612
rect 48924 14572 52920 14600
rect 48924 14560 48930 14572
rect 52914 14560 52920 14572
rect 52972 14560 52978 14612
rect 53469 14603 53527 14609
rect 53469 14569 53481 14603
rect 53515 14600 53527 14603
rect 54113 14603 54171 14609
rect 54113 14600 54125 14603
rect 53515 14572 54125 14600
rect 53515 14569 53527 14572
rect 53469 14563 53527 14569
rect 54113 14569 54125 14572
rect 54159 14569 54171 14603
rect 56870 14600 56876 14612
rect 54113 14563 54171 14569
rect 56428 14572 56876 14600
rect 42518 14492 42524 14544
rect 42576 14532 42582 14544
rect 43809 14535 43867 14541
rect 42576 14504 42659 14532
rect 42576 14492 42582 14504
rect 42631 14473 42659 14504
rect 43809 14501 43821 14535
rect 43855 14532 43867 14535
rect 43990 14532 43996 14544
rect 43855 14504 43996 14532
rect 43855 14501 43867 14504
rect 43809 14495 43867 14501
rect 43990 14492 43996 14504
rect 44048 14492 44054 14544
rect 44174 14492 44180 14544
rect 44232 14532 44238 14544
rect 44361 14535 44419 14541
rect 44361 14532 44373 14535
rect 44232 14504 44373 14532
rect 44232 14492 44238 14504
rect 44361 14501 44373 14504
rect 44407 14501 44419 14535
rect 45370 14532 45376 14544
rect 45331 14504 45376 14532
rect 44361 14495 44419 14501
rect 45370 14492 45376 14504
rect 45428 14492 45434 14544
rect 45830 14492 45836 14544
rect 45888 14532 45894 14544
rect 45888 14504 48176 14532
rect 45888 14492 45894 14504
rect 39117 14467 39175 14473
rect 39117 14433 39129 14467
rect 39163 14433 39175 14467
rect 42613 14467 42671 14473
rect 39117 14427 39175 14433
rect 41616 14436 42564 14464
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14365 20499 14399
rect 20441 14359 20499 14365
rect 20806 14356 20812 14408
rect 20864 14396 20870 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20864 14368 21097 14396
rect 20864 14356 20870 14368
rect 21085 14365 21097 14368
rect 21131 14396 21143 14399
rect 21266 14396 21272 14408
rect 21131 14368 21272 14396
rect 21131 14365 21143 14368
rect 21085 14359 21143 14365
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 22002 14356 22008 14408
rect 22060 14396 22066 14408
rect 22097 14399 22155 14405
rect 22097 14396 22109 14399
rect 22060 14368 22109 14396
rect 22060 14356 22066 14368
rect 22097 14365 22109 14368
rect 22143 14365 22155 14399
rect 22097 14359 22155 14365
rect 23474 14356 23480 14408
rect 23532 14356 23538 14408
rect 26786 14396 26792 14408
rect 26747 14368 26792 14396
rect 26786 14356 26792 14368
rect 26844 14356 26850 14408
rect 27430 14396 27436 14408
rect 27391 14368 27436 14396
rect 27430 14356 27436 14368
rect 27488 14356 27494 14408
rect 27614 14396 27620 14408
rect 27575 14368 27620 14396
rect 27614 14356 27620 14368
rect 27672 14356 27678 14408
rect 29730 14356 29736 14408
rect 29788 14396 29794 14408
rect 29825 14399 29883 14405
rect 29825 14396 29837 14399
rect 29788 14368 29837 14396
rect 29788 14356 29794 14368
rect 29825 14365 29837 14368
rect 29871 14365 29883 14399
rect 37642 14396 37648 14408
rect 29825 14359 29883 14365
rect 37003 14368 37648 14396
rect 20162 14328 20168 14340
rect 19352 14300 20168 14328
rect 20162 14288 20168 14300
rect 20220 14288 20226 14340
rect 20254 14288 20260 14340
rect 20312 14328 20318 14340
rect 21910 14328 21916 14340
rect 20312 14300 21916 14328
rect 20312 14288 20318 14300
rect 21910 14288 21916 14300
rect 21968 14288 21974 14340
rect 22370 14328 22376 14340
rect 22331 14300 22376 14328
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 25406 14288 25412 14340
rect 25464 14288 25470 14340
rect 30101 14331 30159 14337
rect 30101 14297 30113 14331
rect 30147 14328 30159 14331
rect 30837 14331 30895 14337
rect 30837 14328 30849 14331
rect 30147 14300 30849 14328
rect 30147 14297 30159 14300
rect 30101 14291 30159 14297
rect 30837 14297 30849 14300
rect 30883 14297 30895 14331
rect 32214 14328 32220 14340
rect 32062 14300 32220 14328
rect 30837 14291 30895 14297
rect 32214 14288 32220 14300
rect 32272 14288 32278 14340
rect 36538 14328 36544 14340
rect 36202 14300 36544 14328
rect 36538 14288 36544 14300
rect 36596 14288 36602 14340
rect 12342 14260 12348 14272
rect 10652 14232 12348 14260
rect 10652 14220 10658 14232
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 14366 14220 14372 14272
rect 14424 14260 14430 14272
rect 17773 14263 17831 14269
rect 17773 14260 17785 14263
rect 14424 14232 17785 14260
rect 14424 14220 14430 14232
rect 17773 14229 17785 14232
rect 17819 14229 17831 14263
rect 17773 14223 17831 14229
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 21358 14260 21364 14272
rect 18564 14232 21364 14260
rect 18564 14220 18570 14232
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 21453 14263 21511 14269
rect 21453 14229 21465 14263
rect 21499 14260 21511 14263
rect 22186 14260 22192 14272
rect 21499 14232 22192 14260
rect 21499 14229 21511 14232
rect 21453 14223 21511 14229
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 23014 14220 23020 14272
rect 23072 14260 23078 14272
rect 23845 14263 23903 14269
rect 23845 14260 23857 14263
rect 23072 14232 23857 14260
rect 23072 14220 23078 14232
rect 23845 14229 23857 14232
rect 23891 14229 23903 14263
rect 26694 14260 26700 14272
rect 26655 14232 26700 14260
rect 23845 14223 23903 14229
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 28442 14260 28448 14272
rect 28403 14232 28448 14260
rect 28442 14220 28448 14232
rect 28500 14220 28506 14272
rect 32309 14263 32367 14269
rect 32309 14229 32321 14263
rect 32355 14260 32367 14263
rect 32582 14260 32588 14272
rect 32355 14232 32588 14260
rect 32355 14229 32367 14232
rect 32309 14223 32367 14229
rect 32582 14220 32588 14232
rect 32640 14220 32646 14272
rect 35161 14263 35219 14269
rect 35161 14229 35173 14263
rect 35207 14260 35219 14263
rect 37003 14260 37031 14368
rect 37642 14356 37648 14368
rect 37700 14396 37706 14408
rect 38105 14399 38163 14405
rect 38105 14396 38117 14399
rect 37700 14368 38117 14396
rect 37700 14356 37706 14368
rect 38105 14365 38117 14368
rect 38151 14365 38163 14399
rect 38286 14396 38292 14408
rect 38247 14368 38292 14396
rect 38105 14359 38163 14365
rect 38286 14356 38292 14368
rect 38344 14356 38350 14408
rect 40313 14399 40371 14405
rect 40313 14365 40325 14399
rect 40359 14396 40371 14399
rect 40586 14396 40592 14408
rect 40359 14368 40592 14396
rect 40359 14365 40371 14368
rect 40313 14359 40371 14365
rect 40586 14356 40592 14368
rect 40644 14356 40650 14408
rect 40678 14356 40684 14408
rect 40736 14396 40742 14408
rect 40957 14399 41015 14405
rect 40957 14396 40969 14399
rect 40736 14368 40969 14396
rect 40736 14356 40742 14368
rect 40957 14365 40969 14368
rect 41003 14365 41015 14399
rect 40957 14359 41015 14365
rect 41138 14356 41144 14408
rect 41196 14396 41202 14408
rect 41233 14399 41291 14405
rect 41233 14396 41245 14399
rect 41196 14368 41245 14396
rect 41196 14356 41202 14368
rect 41233 14365 41245 14368
rect 41279 14396 41291 14399
rect 41414 14396 41420 14408
rect 41279 14368 41420 14396
rect 41279 14365 41291 14368
rect 41233 14359 41291 14365
rect 41414 14356 41420 14368
rect 41472 14356 41478 14408
rect 39298 14288 39304 14340
rect 39356 14328 39362 14340
rect 41616 14328 41644 14436
rect 41690 14356 41696 14408
rect 41748 14396 41754 14408
rect 41877 14399 41935 14405
rect 41877 14396 41889 14399
rect 41748 14368 41889 14396
rect 41748 14356 41754 14368
rect 41877 14365 41889 14368
rect 41923 14365 41935 14399
rect 42536 14398 42564 14436
rect 42613 14433 42625 14467
rect 42659 14433 42671 14467
rect 42613 14427 42671 14433
rect 44910 14424 44916 14476
rect 44968 14464 44974 14476
rect 45005 14467 45063 14473
rect 45005 14464 45017 14467
rect 44968 14436 45017 14464
rect 44968 14424 44974 14436
rect 45005 14433 45017 14436
rect 45051 14433 45063 14467
rect 46198 14464 46204 14476
rect 46159 14436 46204 14464
rect 45005 14427 45063 14433
rect 46198 14424 46204 14436
rect 46256 14424 46262 14476
rect 46290 14424 46296 14476
rect 46348 14464 46354 14476
rect 46753 14467 46811 14473
rect 46753 14464 46765 14467
rect 46348 14436 46765 14464
rect 46348 14424 46354 14436
rect 46753 14433 46765 14436
rect 46799 14433 46811 14467
rect 46753 14427 46811 14433
rect 48148 14464 48176 14504
rect 48958 14492 48964 14544
rect 49016 14532 49022 14544
rect 49053 14535 49111 14541
rect 49053 14532 49065 14535
rect 49016 14504 49065 14532
rect 49016 14492 49022 14504
rect 49053 14501 49065 14504
rect 49099 14501 49111 14535
rect 49053 14495 49111 14501
rect 51077 14535 51135 14541
rect 51077 14501 51089 14535
rect 51123 14532 51135 14535
rect 51123 14504 52040 14532
rect 51123 14501 51135 14504
rect 51077 14495 51135 14501
rect 50890 14464 50896 14476
rect 48148 14436 50896 14464
rect 42536 14370 42656 14398
rect 42886 14396 42892 14408
rect 41877 14359 41935 14365
rect 39356 14300 41644 14328
rect 39356 14288 39362 14300
rect 41782 14288 41788 14340
rect 41840 14328 41846 14340
rect 42518 14328 42524 14340
rect 41840 14300 42524 14328
rect 41840 14288 41846 14300
rect 42518 14288 42524 14300
rect 42576 14288 42582 14340
rect 42628 14328 42656 14370
rect 42847 14368 42892 14396
rect 42886 14356 42892 14368
rect 42944 14356 42950 14408
rect 43530 14396 43536 14408
rect 43491 14368 43536 14396
rect 43530 14356 43536 14368
rect 43588 14356 43594 14408
rect 44453 14399 44511 14405
rect 44453 14365 44465 14399
rect 44499 14396 44511 14399
rect 44634 14396 44640 14408
rect 44499 14368 44640 14396
rect 44499 14365 44511 14368
rect 44453 14359 44511 14365
rect 44634 14356 44640 14368
rect 44692 14356 44698 14408
rect 45554 14356 45560 14408
rect 45612 14396 45618 14408
rect 45925 14399 45983 14405
rect 45925 14396 45937 14399
rect 45612 14368 45937 14396
rect 45612 14356 45618 14368
rect 45925 14365 45937 14368
rect 45971 14365 45983 14399
rect 45925 14359 45983 14365
rect 46017 14399 46075 14405
rect 46017 14365 46029 14399
rect 46063 14396 46075 14399
rect 46658 14396 46664 14408
rect 46063 14368 46664 14396
rect 46063 14365 46075 14368
rect 46017 14359 46075 14365
rect 46658 14356 46664 14368
rect 46716 14356 46722 14408
rect 46842 14396 46848 14408
rect 46803 14368 46848 14396
rect 46842 14356 46848 14368
rect 46900 14356 46906 14408
rect 48148 14396 48176 14436
rect 50890 14424 50896 14436
rect 50948 14424 50954 14476
rect 51813 14467 51871 14473
rect 51813 14433 51825 14467
rect 51859 14464 51871 14467
rect 51902 14464 51908 14476
rect 51859 14436 51908 14464
rect 51859 14433 51871 14436
rect 51813 14427 51871 14433
rect 51902 14424 51908 14436
rect 51960 14424 51966 14476
rect 52012 14464 52040 14504
rect 52362 14492 52368 14544
rect 52420 14532 52426 14544
rect 52420 14504 54340 14532
rect 52420 14492 52426 14504
rect 52012 14436 53052 14464
rect 48225 14399 48283 14405
rect 48225 14396 48237 14399
rect 48148 14368 48237 14396
rect 48225 14365 48237 14368
rect 48271 14365 48283 14399
rect 48225 14359 48283 14365
rect 48314 14356 48320 14408
rect 48372 14396 48378 14408
rect 48958 14396 48964 14408
rect 48372 14368 48417 14396
rect 48919 14368 48964 14396
rect 48372 14356 48378 14368
rect 48958 14356 48964 14368
rect 49016 14356 49022 14408
rect 49142 14396 49148 14408
rect 49103 14368 49148 14396
rect 49142 14356 49148 14368
rect 49200 14356 49206 14408
rect 50709 14399 50767 14405
rect 50709 14365 50721 14399
rect 50755 14396 50767 14399
rect 51350 14396 51356 14408
rect 50755 14368 51356 14396
rect 50755 14365 50767 14368
rect 50709 14359 50767 14365
rect 51350 14356 51356 14368
rect 51408 14356 51414 14408
rect 51442 14356 51448 14408
rect 51500 14396 51506 14408
rect 51721 14399 51779 14405
rect 51721 14396 51733 14399
rect 51500 14368 51733 14396
rect 51500 14356 51506 14368
rect 51721 14365 51733 14368
rect 51767 14396 51779 14399
rect 51767 14368 52776 14396
rect 51767 14365 51779 14368
rect 51721 14359 51779 14365
rect 44818 14328 44824 14340
rect 42628 14300 44824 14328
rect 44818 14288 44824 14300
rect 44876 14288 44882 14340
rect 45186 14288 45192 14340
rect 45244 14328 45250 14340
rect 45830 14328 45836 14340
rect 45244 14300 45836 14328
rect 45244 14288 45250 14300
rect 45830 14288 45836 14300
rect 45888 14328 45894 14340
rect 48501 14331 48559 14337
rect 45888 14300 48176 14328
rect 45888 14288 45894 14300
rect 35207 14232 37031 14260
rect 35207 14229 35219 14232
rect 35161 14223 35219 14229
rect 37090 14220 37096 14272
rect 37148 14260 37154 14272
rect 37553 14263 37611 14269
rect 37553 14260 37565 14263
rect 37148 14232 37565 14260
rect 37148 14220 37154 14232
rect 37553 14229 37565 14232
rect 37599 14260 37611 14263
rect 40126 14260 40132 14272
rect 37599 14232 40132 14260
rect 37599 14229 37611 14232
rect 37553 14223 37611 14229
rect 40126 14220 40132 14232
rect 40184 14220 40190 14272
rect 40405 14263 40463 14269
rect 40405 14229 40417 14263
rect 40451 14260 40463 14263
rect 42058 14260 42064 14272
rect 40451 14232 42064 14260
rect 40451 14229 40463 14232
rect 40405 14223 40463 14229
rect 42058 14220 42064 14232
rect 42116 14220 42122 14272
rect 42153 14263 42211 14269
rect 42153 14229 42165 14263
rect 42199 14260 42211 14263
rect 42978 14260 42984 14272
rect 42199 14232 42984 14260
rect 42199 14229 42211 14232
rect 42153 14223 42211 14229
rect 42978 14220 42984 14232
rect 43036 14260 43042 14272
rect 43990 14260 43996 14272
rect 43036 14232 43996 14260
rect 43036 14220 43042 14232
rect 43990 14220 43996 14232
rect 44048 14220 44054 14272
rect 45465 14263 45523 14269
rect 45465 14229 45477 14263
rect 45511 14260 45523 14263
rect 45922 14260 45928 14272
rect 45511 14232 45928 14260
rect 45511 14229 45523 14232
rect 45465 14223 45523 14229
rect 45922 14220 45928 14232
rect 45980 14220 45986 14272
rect 47210 14260 47216 14272
rect 47171 14232 47216 14260
rect 47210 14220 47216 14232
rect 47268 14220 47274 14272
rect 47486 14220 47492 14272
rect 47544 14260 47550 14272
rect 48041 14263 48099 14269
rect 48041 14260 48053 14263
rect 47544 14232 48053 14260
rect 47544 14220 47550 14232
rect 48041 14229 48053 14232
rect 48087 14229 48099 14263
rect 48148 14260 48176 14300
rect 48501 14297 48513 14331
rect 48547 14328 48559 14331
rect 51166 14328 51172 14340
rect 48547 14300 51172 14328
rect 48547 14297 48559 14300
rect 48501 14291 48559 14297
rect 51166 14288 51172 14300
rect 51224 14288 51230 14340
rect 52748 14337 52776 14368
rect 52549 14331 52607 14337
rect 52549 14328 52561 14331
rect 51828 14300 52561 14328
rect 48958 14260 48964 14272
rect 48148 14232 48964 14260
rect 48041 14223 48099 14229
rect 48958 14220 48964 14232
rect 49016 14220 49022 14272
rect 50338 14220 50344 14272
rect 50396 14260 50402 14272
rect 50525 14263 50583 14269
rect 50525 14260 50537 14263
rect 50396 14232 50537 14260
rect 50396 14220 50402 14232
rect 50525 14229 50537 14232
rect 50571 14229 50583 14263
rect 50525 14223 50583 14229
rect 50706 14220 50712 14272
rect 50764 14260 50770 14272
rect 50801 14263 50859 14269
rect 50801 14260 50813 14263
rect 50764 14232 50813 14260
rect 50764 14220 50770 14232
rect 50801 14229 50813 14232
rect 50847 14229 50859 14263
rect 50801 14223 50859 14229
rect 50890 14220 50896 14272
rect 50948 14260 50954 14272
rect 51828 14260 51856 14300
rect 52549 14297 52561 14300
rect 52595 14297 52607 14331
rect 52549 14291 52607 14297
rect 52733 14331 52791 14337
rect 52733 14297 52745 14331
rect 52779 14328 52791 14331
rect 52914 14328 52920 14340
rect 52779 14300 52920 14328
rect 52779 14297 52791 14300
rect 52733 14291 52791 14297
rect 52914 14288 52920 14300
rect 52972 14288 52978 14340
rect 53024 14328 53052 14436
rect 53190 14424 53196 14476
rect 53248 14464 53254 14476
rect 54312 14473 54340 14504
rect 53561 14467 53619 14473
rect 53561 14464 53573 14467
rect 53248 14436 53573 14464
rect 53248 14424 53254 14436
rect 53561 14433 53573 14436
rect 53607 14433 53619 14467
rect 53561 14427 53619 14433
rect 54297 14467 54355 14473
rect 54297 14433 54309 14467
rect 54343 14433 54355 14467
rect 54297 14427 54355 14433
rect 53282 14396 53288 14408
rect 53243 14368 53288 14396
rect 53282 14356 53288 14368
rect 53340 14356 53346 14408
rect 53374 14356 53380 14408
rect 53432 14396 53438 14408
rect 53432 14368 53477 14396
rect 53432 14356 53438 14368
rect 53650 14356 53656 14408
rect 53708 14396 53714 14408
rect 54018 14396 54024 14408
rect 53708 14368 54024 14396
rect 53708 14356 53714 14368
rect 54018 14356 54024 14368
rect 54076 14356 54082 14408
rect 54478 14356 54484 14408
rect 54536 14396 54542 14408
rect 56428 14405 56456 14572
rect 56870 14560 56876 14572
rect 56928 14560 56934 14612
rect 57146 14560 57152 14612
rect 57204 14600 57210 14612
rect 58161 14603 58219 14609
rect 58161 14600 58173 14603
rect 57204 14572 58173 14600
rect 57204 14560 57210 14572
rect 58161 14569 58173 14572
rect 58207 14569 58219 14603
rect 58161 14563 58219 14569
rect 56686 14464 56692 14476
rect 56647 14436 56692 14464
rect 56686 14424 56692 14436
rect 56744 14424 56750 14476
rect 56413 14399 56471 14405
rect 56413 14396 56425 14399
rect 54536 14368 56425 14396
rect 54536 14356 54542 14368
rect 56413 14365 56425 14368
rect 56459 14365 56471 14399
rect 56413 14359 56471 14365
rect 53466 14328 53472 14340
rect 53024 14300 53472 14328
rect 53466 14288 53472 14300
rect 53524 14288 53530 14340
rect 57330 14288 57336 14340
rect 57388 14288 57394 14340
rect 50948 14232 51856 14260
rect 50948 14220 50954 14232
rect 51902 14220 51908 14272
rect 51960 14260 51966 14272
rect 52089 14263 52147 14269
rect 52089 14260 52101 14263
rect 51960 14232 52101 14260
rect 51960 14220 51966 14232
rect 52089 14229 52101 14232
rect 52135 14229 52147 14263
rect 52089 14223 52147 14229
rect 54297 14263 54355 14269
rect 54297 14229 54309 14263
rect 54343 14260 54355 14263
rect 56134 14260 56140 14272
rect 54343 14232 56140 14260
rect 54343 14229 54355 14232
rect 54297 14223 54355 14229
rect 56134 14220 56140 14232
rect 56192 14220 56198 14272
rect 1104 14170 58880 14192
rect 1104 14118 15398 14170
rect 15450 14118 15462 14170
rect 15514 14118 15526 14170
rect 15578 14118 15590 14170
rect 15642 14118 15654 14170
rect 15706 14118 29846 14170
rect 29898 14118 29910 14170
rect 29962 14118 29974 14170
rect 30026 14118 30038 14170
rect 30090 14118 30102 14170
rect 30154 14118 44294 14170
rect 44346 14118 44358 14170
rect 44410 14118 44422 14170
rect 44474 14118 44486 14170
rect 44538 14118 44550 14170
rect 44602 14118 58880 14170
rect 1104 14096 58880 14118
rect 6822 14056 6828 14068
rect 6783 14028 6828 14056
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 11422 14056 11428 14068
rect 7944 14028 11428 14056
rect 7944 13932 7972 14028
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 11532 14028 11744 14056
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 8076 13960 9522 13988
rect 8076 13948 8082 13960
rect 10410 13948 10416 14000
rect 10468 13988 10474 14000
rect 11532 13988 11560 14028
rect 10468 13960 11560 13988
rect 11716 13988 11744 14028
rect 11790 14016 11796 14068
rect 11848 14056 11854 14068
rect 12253 14059 12311 14065
rect 12253 14056 12265 14059
rect 11848 14028 12265 14056
rect 11848 14016 11854 14028
rect 12253 14025 12265 14028
rect 12299 14025 12311 14059
rect 12253 14019 12311 14025
rect 12342 14016 12348 14068
rect 12400 14056 12406 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12400 14028 12909 14056
rect 12400 14016 12406 14028
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 16022 14056 16028 14068
rect 12897 14019 12955 14025
rect 13096 14028 16028 14056
rect 11716 13960 12480 13988
rect 10468 13948 10474 13960
rect 6730 13920 6736 13932
rect 6691 13892 6736 13920
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 7926 13920 7932 13932
rect 7839 13892 7932 13920
rect 7926 13880 7932 13892
rect 7984 13880 7990 13932
rect 8754 13920 8760 13932
rect 8715 13892 8760 13920
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13920 11851 13923
rect 12342 13920 12348 13932
rect 11839 13892 12348 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 12452 13929 12480 13960
rect 13096 13929 13124 14028
rect 16022 14016 16028 14028
rect 16080 14016 16086 14068
rect 16117 14059 16175 14065
rect 16117 14025 16129 14059
rect 16163 14056 16175 14059
rect 17126 14056 17132 14068
rect 16163 14028 17132 14056
rect 16163 14025 16175 14028
rect 16117 14019 16175 14025
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 17310 14056 17316 14068
rect 17271 14028 17316 14056
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 18506 14056 18512 14068
rect 18467 14028 18512 14056
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 22830 14056 22836 14068
rect 18616 14028 22836 14056
rect 17954 13988 17960 14000
rect 15870 13960 17960 13988
rect 17954 13948 17960 13960
rect 18012 13948 18018 14000
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13817 13923 13875 13929
rect 13817 13889 13829 13923
rect 13863 13920 13875 13923
rect 13998 13920 14004 13932
rect 13863 13892 14004 13920
rect 13863 13889 13875 13892
rect 13817 13883 13875 13889
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 16574 13880 16580 13932
rect 16632 13920 16638 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16632 13892 16681 13920
rect 16632 13880 16638 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 17405 13923 17463 13929
rect 17405 13889 17417 13923
rect 17451 13889 17463 13923
rect 17405 13883 17463 13889
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18524 13920 18552 14016
rect 18095 13892 18552 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 8018 13852 8024 13864
rect 7979 13824 8024 13852
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 9214 13852 9220 13864
rect 9175 13824 9220 13852
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 10965 13855 11023 13861
rect 10965 13852 10977 13855
rect 10744 13824 10977 13852
rect 10744 13812 10750 13824
rect 10965 13821 10977 13824
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 11701 13855 11759 13861
rect 11701 13821 11713 13855
rect 11747 13852 11759 13855
rect 13906 13852 13912 13864
rect 11747 13824 13912 13852
rect 11747 13821 11759 13824
rect 11701 13815 11759 13821
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14734 13852 14740 13864
rect 14415 13824 14740 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 17420 13852 17448 13883
rect 18616 13852 18644 14028
rect 22830 14016 22836 14028
rect 22888 14016 22894 14068
rect 23934 14056 23940 14068
rect 23895 14028 23940 14056
rect 23934 14016 23940 14028
rect 23992 14056 23998 14068
rect 27430 14056 27436 14068
rect 23992 14028 27436 14056
rect 23992 14016 23998 14028
rect 27430 14016 27436 14028
rect 27488 14016 27494 14068
rect 29549 14059 29607 14065
rect 29549 14025 29561 14059
rect 29595 14056 29607 14059
rect 29730 14056 29736 14068
rect 29595 14028 29736 14056
rect 29595 14025 29607 14028
rect 29549 14019 29607 14025
rect 29730 14016 29736 14028
rect 29788 14056 29794 14068
rect 33229 14059 33287 14065
rect 29788 14028 31754 14056
rect 29788 14016 29794 14028
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 21177 13991 21235 13997
rect 18748 13960 18814 13988
rect 18748 13948 18754 13960
rect 21177 13957 21189 13991
rect 21223 13988 21235 13991
rect 22465 13991 22523 13997
rect 22465 13988 22477 13991
rect 21223 13960 22477 13988
rect 21223 13957 21235 13960
rect 21177 13951 21235 13957
rect 22465 13957 22477 13960
rect 22511 13957 22523 13991
rect 24394 13988 24400 14000
rect 23690 13960 24400 13988
rect 22465 13951 22523 13957
rect 24394 13948 24400 13960
rect 24452 13948 24458 14000
rect 26694 13988 26700 14000
rect 25898 13960 26700 13988
rect 26694 13948 26700 13960
rect 26752 13948 26758 14000
rect 29638 13988 29644 14000
rect 29302 13960 29644 13988
rect 29638 13948 29644 13960
rect 29696 13948 29702 14000
rect 30561 13991 30619 13997
rect 30561 13957 30573 13991
rect 30607 13988 30619 13991
rect 30607 13960 31156 13988
rect 30607 13957 30619 13960
rect 30561 13951 30619 13957
rect 20254 13880 20260 13932
rect 20312 13920 20318 13932
rect 20312 13892 20357 13920
rect 20312 13880 20318 13892
rect 20990 13880 20996 13932
rect 21048 13920 21054 13932
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 21048 13892 21097 13920
rect 21048 13880 21054 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 26973 13923 27031 13929
rect 26973 13920 26985 13923
rect 26292 13892 26985 13920
rect 26292 13880 26298 13892
rect 26973 13889 26985 13892
rect 27019 13889 27031 13923
rect 27798 13920 27804 13932
rect 27759 13892 27804 13920
rect 26973 13883 27031 13889
rect 27798 13880 27804 13892
rect 27856 13880 27862 13932
rect 30285 13923 30343 13929
rect 30285 13889 30297 13923
rect 30331 13920 30343 13923
rect 31018 13920 31024 13932
rect 30331 13892 31024 13920
rect 30331 13889 30343 13892
rect 30285 13883 30343 13889
rect 31018 13880 31024 13892
rect 31076 13880 31082 13932
rect 19978 13852 19984 13864
rect 17420 13824 18644 13852
rect 18708 13824 19984 13852
rect 7834 13744 7840 13796
rect 7892 13784 7898 13796
rect 7892 13756 9352 13784
rect 7892 13744 7898 13756
rect 9324 13716 9352 13756
rect 11422 13744 11428 13796
rect 11480 13784 11486 13796
rect 13538 13784 13544 13796
rect 11480 13756 13544 13784
rect 11480 13744 11486 13756
rect 13538 13744 13544 13756
rect 13596 13784 13602 13796
rect 13633 13787 13691 13793
rect 13633 13784 13645 13787
rect 13596 13756 13645 13784
rect 13596 13744 13602 13756
rect 13633 13753 13645 13756
rect 13679 13753 13691 13787
rect 13633 13747 13691 13753
rect 17957 13787 18015 13793
rect 17957 13753 17969 13787
rect 18003 13784 18015 13787
rect 18708 13784 18736 13824
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 22189 13855 22247 13861
rect 22189 13821 22201 13855
rect 22235 13852 22247 13855
rect 23198 13852 23204 13864
rect 22235 13824 23204 13852
rect 22235 13821 22247 13824
rect 22189 13815 22247 13821
rect 23198 13812 23204 13824
rect 23256 13812 23262 13864
rect 24118 13812 24124 13864
rect 24176 13852 24182 13864
rect 24397 13855 24455 13861
rect 24397 13852 24409 13855
rect 24176 13824 24409 13852
rect 24176 13812 24182 13824
rect 24397 13821 24409 13824
rect 24443 13852 24455 13855
rect 24762 13852 24768 13864
rect 24443 13824 24768 13852
rect 24443 13821 24455 13824
rect 24397 13815 24455 13821
rect 24762 13812 24768 13824
rect 24820 13812 24826 13864
rect 26145 13855 26203 13861
rect 26145 13821 26157 13855
rect 26191 13852 26203 13855
rect 27062 13852 27068 13864
rect 26191 13824 26924 13852
rect 27023 13824 27068 13852
rect 26191 13821 26203 13824
rect 26145 13815 26203 13821
rect 18003 13756 18736 13784
rect 26896 13784 26924 13824
rect 27062 13812 27068 13824
rect 27120 13812 27126 13864
rect 27522 13852 27528 13864
rect 27172 13824 27528 13852
rect 27172 13784 27200 13824
rect 27522 13812 27528 13824
rect 27580 13812 27586 13864
rect 28074 13852 28080 13864
rect 28035 13824 28080 13852
rect 28074 13812 28080 13824
rect 28132 13812 28138 13864
rect 30561 13855 30619 13861
rect 30561 13821 30573 13855
rect 30607 13852 30619 13855
rect 30742 13852 30748 13864
rect 30607 13824 30748 13852
rect 30607 13821 30619 13824
rect 30561 13815 30619 13821
rect 30742 13812 30748 13824
rect 30800 13812 30806 13864
rect 31128 13861 31156 13960
rect 31202 13880 31208 13932
rect 31260 13920 31266 13932
rect 31726 13920 31754 14028
rect 33229 14025 33241 14059
rect 33275 14056 33287 14059
rect 33275 14028 37780 14056
rect 33275 14025 33287 14028
rect 33229 14019 33287 14025
rect 34238 13988 34244 14000
rect 32600 13960 34244 13988
rect 32401 13923 32459 13929
rect 32401 13920 32413 13923
rect 31260 13892 31305 13920
rect 31726 13892 32413 13920
rect 31260 13880 31266 13892
rect 32401 13889 32413 13892
rect 32447 13889 32459 13923
rect 32401 13883 32459 13889
rect 31113 13855 31171 13861
rect 31113 13821 31125 13855
rect 31159 13821 31171 13855
rect 31113 13815 31171 13821
rect 31294 13812 31300 13864
rect 31352 13852 31358 13864
rect 32600 13852 32628 13960
rect 34238 13948 34244 13960
rect 34296 13948 34302 14000
rect 34882 13948 34888 14000
rect 34940 13948 34946 14000
rect 37752 13997 37780 14028
rect 41690 14016 41696 14068
rect 41748 14056 41754 14068
rect 43625 14059 43683 14065
rect 41748 14028 43392 14056
rect 41748 14016 41754 14028
rect 37737 13991 37795 13997
rect 37737 13957 37749 13991
rect 37783 13957 37795 13991
rect 37737 13951 37795 13957
rect 40678 13948 40684 14000
rect 40736 13988 40742 14000
rect 40736 13960 42472 13988
rect 40736 13948 40742 13960
rect 33594 13880 33600 13932
rect 33652 13920 33658 13932
rect 33873 13923 33931 13929
rect 33873 13920 33885 13923
rect 33652 13892 33885 13920
rect 33652 13880 33658 13892
rect 33873 13889 33885 13892
rect 33919 13889 33931 13923
rect 40034 13920 40040 13932
rect 39995 13892 40040 13920
rect 33873 13883 33931 13889
rect 40034 13880 40040 13892
rect 40092 13880 40098 13932
rect 40954 13920 40960 13932
rect 40915 13892 40960 13920
rect 40954 13880 40960 13892
rect 41012 13880 41018 13932
rect 41690 13920 41696 13932
rect 41651 13892 41696 13920
rect 41690 13880 41696 13892
rect 41748 13880 41754 13932
rect 42444 13929 42472 13960
rect 42518 13948 42524 14000
rect 42576 13988 42582 14000
rect 42576 13960 42840 13988
rect 42576 13948 42582 13960
rect 42429 13923 42487 13929
rect 42429 13889 42441 13923
rect 42475 13889 42487 13923
rect 42702 13920 42708 13932
rect 42663 13892 42708 13920
rect 42429 13883 42487 13889
rect 42702 13880 42708 13892
rect 42760 13880 42766 13932
rect 42812 13920 42840 13960
rect 43364 13929 43392 14028
rect 43625 14025 43637 14059
rect 43671 14056 43683 14059
rect 43990 14056 43996 14068
rect 43671 14028 43996 14056
rect 43671 14025 43683 14028
rect 43625 14019 43683 14025
rect 43990 14016 43996 14028
rect 44048 14016 44054 14068
rect 45005 14059 45063 14065
rect 45005 14025 45017 14059
rect 45051 14056 45063 14059
rect 45462 14056 45468 14068
rect 45051 14028 45468 14056
rect 45051 14025 45063 14028
rect 45005 14019 45063 14025
rect 45462 14016 45468 14028
rect 45520 14016 45526 14068
rect 46109 14059 46167 14065
rect 46109 14025 46121 14059
rect 46155 14056 46167 14059
rect 46290 14056 46296 14068
rect 46155 14028 46296 14056
rect 46155 14025 46167 14028
rect 46109 14019 46167 14025
rect 46290 14016 46296 14028
rect 46348 14016 46354 14068
rect 46658 14056 46664 14068
rect 46619 14028 46664 14056
rect 46658 14016 46664 14028
rect 46716 14016 46722 14068
rect 48038 14056 48044 14068
rect 46768 14028 48044 14056
rect 43438 13948 43444 14000
rect 43496 13988 43502 14000
rect 44818 13988 44824 14000
rect 43496 13960 44680 13988
rect 44779 13960 44824 13988
rect 43496 13948 43502 13960
rect 43349 13923 43407 13929
rect 42812 13892 43300 13920
rect 31352 13824 32628 13852
rect 31352 13812 31358 13824
rect 32674 13812 32680 13864
rect 32732 13852 32738 13864
rect 34149 13855 34207 13861
rect 34149 13852 34161 13855
rect 32732 13824 32777 13852
rect 33980 13824 34161 13852
rect 32732 13812 32738 13824
rect 26896 13756 27200 13784
rect 18003 13753 18015 13756
rect 17957 13747 18015 13753
rect 29086 13744 29092 13796
rect 29144 13784 29150 13796
rect 31573 13787 31631 13793
rect 29144 13756 30512 13784
rect 29144 13744 29150 13756
rect 10701 13719 10759 13725
rect 10701 13716 10713 13719
rect 9324 13688 10713 13716
rect 10701 13685 10713 13688
rect 10747 13685 10759 13719
rect 10701 13679 10759 13685
rect 14632 13719 14690 13725
rect 14632 13685 14644 13719
rect 14678 13716 14690 13719
rect 15838 13716 15844 13728
rect 14678 13688 15844 13716
rect 14678 13685 14690 13688
rect 14632 13679 14690 13685
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 19610 13676 19616 13728
rect 19668 13716 19674 13728
rect 19993 13719 20051 13725
rect 19993 13716 20005 13719
rect 19668 13688 20005 13716
rect 19668 13676 19674 13688
rect 19993 13685 20005 13688
rect 20039 13685 20051 13719
rect 19993 13679 20051 13685
rect 24660 13719 24718 13725
rect 24660 13685 24672 13719
rect 24706 13716 24718 13719
rect 30190 13716 30196 13728
rect 24706 13688 30196 13716
rect 24706 13685 24718 13688
rect 24660 13679 24718 13685
rect 30190 13676 30196 13688
rect 30248 13676 30254 13728
rect 30374 13716 30380 13728
rect 30335 13688 30380 13716
rect 30374 13676 30380 13688
rect 30432 13676 30438 13728
rect 30484 13716 30512 13756
rect 31573 13753 31585 13787
rect 31619 13784 31631 13787
rect 32398 13784 32404 13796
rect 31619 13756 32404 13784
rect 31619 13753 31631 13756
rect 31573 13747 31631 13753
rect 32398 13744 32404 13756
rect 32456 13744 32462 13796
rect 33980 13784 34008 13824
rect 34149 13821 34161 13824
rect 34195 13821 34207 13855
rect 34149 13815 34207 13821
rect 34238 13812 34244 13864
rect 34296 13852 34302 13864
rect 35621 13855 35679 13861
rect 35621 13852 35633 13855
rect 34296 13824 35633 13852
rect 34296 13812 34302 13824
rect 35621 13821 35633 13824
rect 35667 13821 35679 13855
rect 35621 13815 35679 13821
rect 37553 13855 37611 13861
rect 37553 13821 37565 13855
rect 37599 13852 37611 13855
rect 39298 13852 39304 13864
rect 37599 13824 39304 13852
rect 37599 13821 37611 13824
rect 37553 13815 37611 13821
rect 39298 13812 39304 13824
rect 39356 13812 39362 13864
rect 39390 13812 39396 13864
rect 39448 13852 39454 13864
rect 40678 13852 40684 13864
rect 39448 13824 39493 13852
rect 40236 13824 40684 13852
rect 39448 13812 39454 13824
rect 40236 13793 40264 13824
rect 40678 13812 40684 13824
rect 40736 13812 40742 13864
rect 43272 13852 43300 13892
rect 43349 13889 43361 13923
rect 43395 13889 43407 13923
rect 43349 13883 43407 13889
rect 44269 13923 44327 13929
rect 44269 13889 44281 13923
rect 44315 13889 44327 13923
rect 44269 13883 44327 13889
rect 44284 13852 44312 13883
rect 43272 13824 44312 13852
rect 44652 13852 44680 13960
rect 44818 13948 44824 13960
rect 44876 13948 44882 14000
rect 44910 13948 44916 14000
rect 44968 13988 44974 14000
rect 45094 13988 45100 14000
rect 44968 13960 45100 13988
rect 44968 13948 44974 13960
rect 45094 13948 45100 13960
rect 45152 13948 45158 14000
rect 45186 13920 45192 13932
rect 45147 13892 45192 13920
rect 45186 13880 45192 13892
rect 45244 13880 45250 13932
rect 45373 13923 45431 13929
rect 45373 13889 45385 13923
rect 45419 13920 45431 13923
rect 45830 13920 45836 13932
rect 45419 13892 45836 13920
rect 45419 13889 45431 13892
rect 45373 13883 45431 13889
rect 45830 13880 45836 13892
rect 45888 13880 45894 13932
rect 46014 13880 46020 13932
rect 46072 13920 46078 13932
rect 46768 13929 46796 14028
rect 48038 14016 48044 14028
rect 48096 14016 48102 14068
rect 48222 14016 48228 14068
rect 48280 14056 48286 14068
rect 48280 14028 49188 14056
rect 48280 14016 48286 14028
rect 47210 13948 47216 14000
rect 47268 13988 47274 14000
rect 47857 13991 47915 13997
rect 47857 13988 47869 13991
rect 47268 13960 47869 13988
rect 47268 13948 47274 13960
rect 47857 13957 47869 13960
rect 47903 13957 47915 13991
rect 47857 13951 47915 13957
rect 48130 13948 48136 14000
rect 48188 13988 48194 14000
rect 49160 13988 49188 14028
rect 49234 14016 49240 14068
rect 49292 14056 49298 14068
rect 49329 14059 49387 14065
rect 49329 14056 49341 14059
rect 49292 14028 49341 14056
rect 49292 14016 49298 14028
rect 49329 14025 49341 14028
rect 49375 14056 49387 14059
rect 50614 14056 50620 14068
rect 49375 14028 50016 14056
rect 50527 14028 50620 14056
rect 49375 14025 49387 14028
rect 49329 14019 49387 14025
rect 49988 13997 50016 14028
rect 50614 14016 50620 14028
rect 50672 14056 50678 14068
rect 51258 14056 51264 14068
rect 50672 14028 51264 14056
rect 50672 14016 50678 14028
rect 51258 14016 51264 14028
rect 51316 14016 51322 14068
rect 53834 14056 53840 14068
rect 53795 14028 53840 14056
rect 53834 14016 53840 14028
rect 53892 14016 53898 14068
rect 54665 14059 54723 14065
rect 54665 14025 54677 14059
rect 54711 14056 54723 14059
rect 55582 14056 55588 14068
rect 54711 14028 55588 14056
rect 54711 14025 54723 14028
rect 54665 14019 54723 14025
rect 55582 14016 55588 14028
rect 55640 14016 55646 14068
rect 57238 14056 57244 14068
rect 57199 14028 57244 14056
rect 57238 14016 57244 14028
rect 57296 14016 57302 14068
rect 49789 13991 49847 13997
rect 49789 13988 49801 13991
rect 48188 13960 48346 13988
rect 49160 13960 49801 13988
rect 48188 13948 48194 13960
rect 49789 13957 49801 13960
rect 49835 13957 49847 13991
rect 49789 13951 49847 13957
rect 49973 13991 50031 13997
rect 49973 13957 49985 13991
rect 50019 13957 50031 13991
rect 50890 13988 50896 14000
rect 49973 13951 50031 13957
rect 50540 13960 50896 13988
rect 50540 13929 50568 13960
rect 50890 13948 50896 13960
rect 50948 13948 50954 14000
rect 53466 13948 53472 14000
rect 53524 13988 53530 14000
rect 57256 13988 57284 14016
rect 53524 13960 56272 13988
rect 57256 13960 58112 13988
rect 53524 13948 53530 13960
rect 46569 13923 46627 13929
rect 46569 13920 46581 13923
rect 46072 13892 46581 13920
rect 46072 13880 46078 13892
rect 46569 13889 46581 13892
rect 46615 13889 46627 13923
rect 46569 13883 46627 13889
rect 46753 13923 46811 13929
rect 46753 13889 46765 13923
rect 46799 13889 46811 13923
rect 46753 13883 46811 13889
rect 50525 13923 50583 13929
rect 50525 13889 50537 13923
rect 50571 13889 50583 13923
rect 50525 13883 50583 13889
rect 50709 13923 50767 13929
rect 50709 13889 50721 13923
rect 50755 13920 50767 13923
rect 51166 13920 51172 13932
rect 50755 13892 51172 13920
rect 50755 13889 50767 13892
rect 50709 13883 50767 13889
rect 51166 13880 51172 13892
rect 51224 13920 51230 13932
rect 52178 13920 52184 13932
rect 51224 13892 52184 13920
rect 51224 13880 51230 13892
rect 52178 13880 52184 13892
rect 52236 13880 52242 13932
rect 53190 13920 53196 13932
rect 53151 13892 53196 13920
rect 53190 13880 53196 13892
rect 53248 13880 53254 13932
rect 53852 13929 53880 13960
rect 53837 13923 53895 13929
rect 53837 13889 53849 13923
rect 53883 13889 53895 13923
rect 53837 13883 53895 13889
rect 54018 13880 54024 13932
rect 54076 13920 54082 13932
rect 54076 13892 54121 13920
rect 54076 13880 54082 13892
rect 54202 13880 54208 13932
rect 54260 13920 54266 13932
rect 54478 13920 54484 13932
rect 54260 13892 54484 13920
rect 54260 13880 54266 13892
rect 54478 13880 54484 13892
rect 54536 13880 54542 13932
rect 56244 13929 56272 13960
rect 56229 13923 56287 13929
rect 56229 13889 56241 13923
rect 56275 13920 56287 13923
rect 57974 13920 57980 13932
rect 56275 13892 57980 13920
rect 56275 13889 56287 13892
rect 56229 13883 56287 13889
rect 57974 13880 57980 13892
rect 58032 13880 58038 13932
rect 58084 13929 58112 13960
rect 58069 13923 58127 13929
rect 58069 13889 58081 13923
rect 58115 13889 58127 13923
rect 58069 13883 58127 13889
rect 46109 13855 46167 13861
rect 46109 13852 46121 13855
rect 44652 13824 46121 13852
rect 46109 13821 46121 13824
rect 46155 13852 46167 13855
rect 46198 13852 46204 13864
rect 46155 13824 46204 13852
rect 46155 13821 46167 13824
rect 46109 13815 46167 13821
rect 46198 13812 46204 13824
rect 46256 13852 46262 13864
rect 47581 13855 47639 13861
rect 46256 13824 47532 13852
rect 46256 13812 46262 13824
rect 32508 13756 34008 13784
rect 40221 13787 40279 13793
rect 32508 13716 32536 13756
rect 40221 13753 40233 13787
rect 40267 13753 40279 13787
rect 40221 13747 40279 13753
rect 43530 13744 43536 13796
rect 43588 13784 43594 13796
rect 44085 13787 44143 13793
rect 44085 13784 44097 13787
rect 43588 13756 44097 13784
rect 43588 13744 43594 13756
rect 44085 13753 44097 13756
rect 44131 13753 44143 13787
rect 45922 13784 45928 13796
rect 45883 13756 45928 13784
rect 44085 13747 44143 13753
rect 45922 13744 45928 13756
rect 45980 13744 45986 13796
rect 30484 13688 32536 13716
rect 41877 13719 41935 13725
rect 41877 13685 41889 13719
rect 41923 13716 41935 13719
rect 42150 13716 42156 13728
rect 41923 13688 42156 13716
rect 41923 13685 41935 13688
rect 41877 13679 41935 13685
rect 42150 13676 42156 13688
rect 42208 13676 42214 13728
rect 47504 13716 47532 13824
rect 47581 13821 47593 13855
rect 47627 13852 47639 13855
rect 49970 13852 49976 13864
rect 47627 13824 49976 13852
rect 47627 13821 47639 13824
rect 47581 13815 47639 13821
rect 49970 13812 49976 13824
rect 50028 13812 50034 13864
rect 51350 13852 51356 13864
rect 51311 13824 51356 13852
rect 51350 13812 51356 13824
rect 51408 13812 51414 13864
rect 51629 13855 51687 13861
rect 51629 13821 51641 13855
rect 51675 13852 51687 13855
rect 53377 13855 53435 13861
rect 51675 13824 53328 13852
rect 51675 13821 51687 13824
rect 51629 13815 51687 13821
rect 53300 13784 53328 13824
rect 53377 13821 53389 13855
rect 53423 13852 53435 13855
rect 56134 13852 56140 13864
rect 53423 13824 54984 13852
rect 56095 13824 56140 13852
rect 53423 13821 53435 13824
rect 53377 13815 53435 13821
rect 54202 13784 54208 13796
rect 53300 13756 54208 13784
rect 54202 13744 54208 13756
rect 54260 13744 54266 13796
rect 54956 13784 54984 13824
rect 56134 13812 56140 13824
rect 56192 13812 56198 13864
rect 56042 13784 56048 13796
rect 54956 13756 56048 13784
rect 56042 13744 56048 13756
rect 56100 13744 56106 13796
rect 49142 13716 49148 13728
rect 47504 13688 49148 13716
rect 49142 13676 49148 13688
rect 49200 13676 49206 13728
rect 56505 13719 56563 13725
rect 56505 13685 56517 13719
rect 56551 13716 56563 13719
rect 56686 13716 56692 13728
rect 56551 13688 56692 13716
rect 56551 13685 56563 13688
rect 56505 13679 56563 13685
rect 56686 13676 56692 13688
rect 56744 13676 56750 13728
rect 57882 13716 57888 13728
rect 57843 13688 57888 13716
rect 57882 13676 57888 13688
rect 57940 13676 57946 13728
rect 1104 13626 58880 13648
rect 1104 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 8302 13626
rect 8354 13574 8366 13626
rect 8418 13574 8430 13626
rect 8482 13574 22622 13626
rect 22674 13574 22686 13626
rect 22738 13574 22750 13626
rect 22802 13574 22814 13626
rect 22866 13574 22878 13626
rect 22930 13574 37070 13626
rect 37122 13574 37134 13626
rect 37186 13574 37198 13626
rect 37250 13574 37262 13626
rect 37314 13574 37326 13626
rect 37378 13574 51518 13626
rect 51570 13574 51582 13626
rect 51634 13574 51646 13626
rect 51698 13574 51710 13626
rect 51762 13574 51774 13626
rect 51826 13574 58880 13626
rect 1104 13552 58880 13574
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 10045 13515 10103 13521
rect 6052 13484 9260 13512
rect 6052 13472 6058 13484
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 7193 13447 7251 13453
rect 7193 13444 7205 13447
rect 6972 13416 7205 13444
rect 6972 13404 6978 13416
rect 7193 13413 7205 13416
rect 7239 13413 7251 13447
rect 9232 13444 9260 13484
rect 10045 13481 10057 13515
rect 10091 13512 10103 13515
rect 10410 13512 10416 13524
rect 10091 13484 10416 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 12253 13515 12311 13521
rect 12253 13481 12265 13515
rect 12299 13512 12311 13515
rect 12434 13512 12440 13524
rect 12299 13484 12440 13512
rect 12299 13481 12311 13484
rect 12253 13475 12311 13481
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 17034 13512 17040 13524
rect 14752 13484 17040 13512
rect 14752 13444 14780 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 20349 13515 20407 13521
rect 20349 13481 20361 13515
rect 20395 13512 20407 13515
rect 24026 13512 24032 13524
rect 20395 13484 24032 13512
rect 20395 13481 20407 13484
rect 20349 13475 20407 13481
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 24394 13472 24400 13524
rect 24452 13512 24458 13524
rect 24489 13515 24547 13521
rect 24489 13512 24501 13515
rect 24452 13484 24501 13512
rect 24452 13472 24458 13484
rect 24489 13481 24501 13484
rect 24535 13481 24547 13515
rect 24489 13475 24547 13481
rect 26786 13472 26792 13524
rect 26844 13512 26850 13524
rect 27341 13515 27399 13521
rect 27341 13512 27353 13515
rect 26844 13484 27353 13512
rect 26844 13472 26850 13484
rect 27341 13481 27353 13484
rect 27387 13481 27399 13515
rect 27341 13475 27399 13481
rect 28074 13472 28080 13524
rect 28132 13512 28138 13524
rect 28721 13515 28779 13521
rect 28721 13512 28733 13515
rect 28132 13484 28733 13512
rect 28132 13472 28138 13484
rect 28721 13481 28733 13484
rect 28767 13481 28779 13515
rect 29638 13512 29644 13524
rect 29599 13484 29644 13512
rect 28721 13475 28779 13481
rect 29638 13472 29644 13484
rect 29696 13472 29702 13524
rect 33962 13512 33968 13524
rect 33923 13484 33968 13512
rect 33962 13472 33968 13484
rect 34020 13472 34026 13524
rect 39301 13515 39359 13521
rect 39301 13481 39313 13515
rect 39347 13512 39359 13515
rect 39942 13512 39948 13524
rect 39347 13484 39948 13512
rect 39347 13481 39359 13484
rect 39301 13475 39359 13481
rect 39942 13472 39948 13484
rect 40000 13472 40006 13524
rect 40034 13472 40040 13524
rect 40092 13512 40098 13524
rect 40313 13515 40371 13521
rect 40313 13512 40325 13515
rect 40092 13484 40325 13512
rect 40092 13472 40098 13484
rect 40313 13481 40325 13484
rect 40359 13512 40371 13515
rect 40586 13512 40592 13524
rect 40359 13484 40592 13512
rect 40359 13481 40371 13484
rect 40313 13475 40371 13481
rect 40586 13472 40592 13484
rect 40644 13512 40650 13524
rect 42610 13512 42616 13524
rect 40644 13484 42616 13512
rect 40644 13472 40650 13484
rect 42610 13472 42616 13484
rect 42668 13472 42674 13524
rect 43809 13515 43867 13521
rect 43809 13481 43821 13515
rect 43855 13512 43867 13515
rect 43990 13512 43996 13524
rect 43855 13484 43996 13512
rect 43855 13481 43867 13484
rect 43809 13475 43867 13481
rect 9232 13416 14780 13444
rect 19337 13447 19395 13453
rect 7193 13407 7251 13413
rect 19337 13413 19349 13447
rect 19383 13444 19395 13447
rect 22370 13444 22376 13456
rect 19383 13416 22376 13444
rect 19383 13413 19395 13416
rect 19337 13407 19395 13413
rect 22370 13404 22376 13416
rect 22428 13404 22434 13456
rect 22462 13404 22468 13456
rect 22520 13444 22526 13456
rect 22520 13416 32720 13444
rect 22520 13404 22526 13416
rect 7653 13379 7711 13385
rect 7653 13345 7665 13379
rect 7699 13376 7711 13379
rect 8018 13376 8024 13388
rect 7699 13348 8024 13376
rect 7699 13345 7711 13348
rect 7653 13339 7711 13345
rect 8018 13336 8024 13348
rect 8076 13336 8082 13388
rect 15286 13376 15292 13388
rect 12406 13348 15292 13376
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 7926 13308 7932 13320
rect 7607 13280 7932 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 11333 13311 11391 13317
rect 11333 13277 11345 13311
rect 11379 13308 11391 13311
rect 12406 13308 12434 13348
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 23845 13379 23903 13385
rect 15804 13348 19288 13376
rect 15804 13336 15810 13348
rect 11379 13280 12434 13308
rect 13541 13311 13599 13317
rect 11379 13277 11391 13280
rect 11333 13271 11391 13277
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 14366 13308 14372 13320
rect 13587 13280 14372 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 19260 13317 19288 13348
rect 23845 13345 23857 13379
rect 23891 13376 23903 13379
rect 24578 13376 24584 13388
rect 23891 13348 24584 13376
rect 23891 13345 23903 13348
rect 23845 13339 23903 13345
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 30561 13379 30619 13385
rect 30561 13345 30573 13379
rect 30607 13376 30619 13379
rect 30742 13376 30748 13388
rect 30607 13348 30748 13376
rect 30607 13345 30619 13348
rect 30561 13339 30619 13345
rect 30742 13336 30748 13348
rect 30800 13336 30806 13388
rect 32582 13376 32588 13388
rect 30944 13348 32588 13376
rect 16853 13311 16911 13317
rect 16853 13308 16865 13311
rect 16080 13280 16125 13308
rect 16776 13280 16865 13308
rect 16080 13268 16086 13280
rect 13906 13200 13912 13252
rect 13964 13240 13970 13252
rect 15749 13243 15807 13249
rect 13964 13212 14582 13240
rect 13964 13200 13970 13212
rect 15749 13209 15761 13243
rect 15795 13240 15807 13243
rect 16574 13240 16580 13252
rect 15795 13212 16580 13240
rect 15795 13209 15807 13212
rect 15749 13203 15807 13209
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8297 13175 8355 13181
rect 8297 13172 8309 13175
rect 8076 13144 8309 13172
rect 8076 13132 8082 13144
rect 8297 13141 8309 13144
rect 8343 13172 8355 13175
rect 9033 13175 9091 13181
rect 9033 13172 9045 13175
rect 8343 13144 9045 13172
rect 8343 13141 8355 13144
rect 8297 13135 8355 13141
rect 9033 13141 9045 13144
rect 9079 13172 9091 13175
rect 13722 13172 13728 13184
rect 9079 13144 13728 13172
rect 9079 13141 9091 13144
rect 9033 13135 9091 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 14274 13172 14280 13184
rect 14235 13144 14280 13172
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 16776 13172 16804 13280
rect 16853 13277 16865 13280
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13308 19303 13311
rect 19886 13308 19892 13320
rect 19291 13280 19892 13308
rect 19291 13277 19303 13280
rect 19245 13271 19303 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 22094 13308 22100 13320
rect 22055 13280 22100 13308
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 24394 13308 24400 13320
rect 24355 13280 24400 13308
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 25593 13311 25651 13317
rect 25593 13277 25605 13311
rect 25639 13308 25651 13311
rect 26234 13308 26240 13320
rect 25639 13280 26240 13308
rect 25639 13277 25651 13280
rect 25593 13271 25651 13277
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 28905 13311 28963 13317
rect 28905 13277 28917 13311
rect 28951 13277 28963 13311
rect 28905 13271 28963 13277
rect 17034 13240 17040 13252
rect 16995 13212 17040 13240
rect 17034 13200 17040 13212
rect 17092 13200 17098 13252
rect 18598 13200 18604 13252
rect 18656 13240 18662 13252
rect 18693 13243 18751 13249
rect 18693 13240 18705 13243
rect 18656 13212 18705 13240
rect 18656 13200 18662 13212
rect 18693 13209 18705 13212
rect 18739 13209 18751 13243
rect 18693 13203 18751 13209
rect 21637 13243 21695 13249
rect 21637 13209 21649 13243
rect 21683 13240 21695 13243
rect 25958 13240 25964 13252
rect 21683 13212 25964 13240
rect 21683 13209 21695 13212
rect 21637 13203 21695 13209
rect 25958 13200 25964 13212
rect 26016 13240 26022 13252
rect 26053 13243 26111 13249
rect 26053 13240 26065 13243
rect 26016 13212 26065 13240
rect 26016 13200 26022 13212
rect 26053 13209 26065 13212
rect 26099 13209 26111 13243
rect 28920 13240 28948 13271
rect 29454 13268 29460 13320
rect 29512 13308 29518 13320
rect 29733 13311 29791 13317
rect 29733 13308 29745 13311
rect 29512 13280 29745 13308
rect 29512 13268 29518 13280
rect 29733 13277 29745 13280
rect 29779 13277 29791 13311
rect 30282 13308 30288 13320
rect 30243 13280 30288 13308
rect 29733 13271 29791 13277
rect 30282 13268 30288 13280
rect 30340 13268 30346 13320
rect 30377 13311 30435 13317
rect 30377 13277 30389 13311
rect 30423 13308 30435 13311
rect 30834 13308 30840 13320
rect 30423 13280 30840 13308
rect 30423 13277 30435 13280
rect 30377 13271 30435 13277
rect 30834 13268 30840 13280
rect 30892 13268 30898 13320
rect 30944 13240 30972 13348
rect 32582 13336 32588 13348
rect 32640 13336 32646 13388
rect 32692 13385 32720 13416
rect 32677 13379 32735 13385
rect 32677 13345 32689 13379
rect 32723 13345 32735 13379
rect 32677 13339 32735 13345
rect 36906 13336 36912 13388
rect 36964 13376 36970 13388
rect 37093 13379 37151 13385
rect 37093 13376 37105 13379
rect 36964 13348 37105 13376
rect 36964 13336 36970 13348
rect 37093 13345 37105 13348
rect 37139 13345 37151 13379
rect 37093 13339 37151 13345
rect 37384 13348 37964 13376
rect 32861 13311 32919 13317
rect 32861 13277 32873 13311
rect 32907 13308 32919 13311
rect 35667 13311 35725 13317
rect 35667 13308 35679 13311
rect 32907 13280 35679 13308
rect 32907 13277 32919 13280
rect 32861 13271 32919 13277
rect 35667 13277 35679 13280
rect 35713 13308 35725 13311
rect 36262 13308 36268 13320
rect 35713 13280 36268 13308
rect 35713 13277 35725 13280
rect 35667 13271 35725 13277
rect 36262 13268 36268 13280
rect 36320 13268 36326 13320
rect 28920 13212 30972 13240
rect 26053 13203 26111 13209
rect 31018 13200 31024 13252
rect 31076 13240 31082 13252
rect 31386 13240 31392 13252
rect 31076 13212 31392 13240
rect 31076 13200 31082 13212
rect 31386 13200 31392 13212
rect 31444 13200 31450 13252
rect 33686 13200 33692 13252
rect 33744 13240 33750 13252
rect 34885 13243 34943 13249
rect 34885 13240 34897 13243
rect 33744 13212 34897 13240
rect 33744 13200 33750 13212
rect 34885 13209 34897 13212
rect 34931 13209 34943 13243
rect 34885 13203 34943 13209
rect 35069 13243 35127 13249
rect 35069 13209 35081 13243
rect 35115 13240 35127 13243
rect 35526 13240 35532 13252
rect 35115 13212 35532 13240
rect 35115 13209 35127 13212
rect 35069 13203 35127 13209
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 35912 13212 36110 13240
rect 18782 13172 18788 13184
rect 16776 13144 18788 13172
rect 18782 13132 18788 13144
rect 18840 13132 18846 13184
rect 25406 13132 25412 13184
rect 25464 13172 25470 13184
rect 25501 13175 25559 13181
rect 25501 13172 25513 13175
rect 25464 13144 25513 13172
rect 25464 13132 25470 13144
rect 25501 13141 25513 13144
rect 25547 13141 25559 13175
rect 25501 13135 25559 13141
rect 30561 13175 30619 13181
rect 30561 13141 30573 13175
rect 30607 13172 30619 13175
rect 32214 13172 32220 13184
rect 30607 13144 32220 13172
rect 30607 13141 30619 13144
rect 30561 13135 30619 13141
rect 32214 13132 32220 13144
rect 32272 13132 32278 13184
rect 33134 13132 33140 13184
rect 33192 13172 33198 13184
rect 33321 13175 33379 13181
rect 33321 13172 33333 13175
rect 33192 13144 33333 13172
rect 33192 13132 33198 13144
rect 33321 13141 33333 13144
rect 33367 13141 33379 13175
rect 33321 13135 33379 13141
rect 34790 13132 34796 13184
rect 34848 13172 34854 13184
rect 35912 13172 35940 13212
rect 37384 13172 37412 13348
rect 37936 13317 37964 13348
rect 40678 13336 40684 13388
rect 40736 13376 40742 13388
rect 40957 13379 41015 13385
rect 40957 13376 40969 13379
rect 40736 13348 40969 13376
rect 40736 13336 40742 13348
rect 40957 13345 40969 13348
rect 41003 13345 41015 13379
rect 42610 13376 42616 13388
rect 42571 13348 42616 13376
rect 40957 13339 41015 13345
rect 42610 13336 42616 13348
rect 42668 13336 42674 13388
rect 37461 13311 37519 13317
rect 37461 13277 37473 13311
rect 37507 13277 37519 13311
rect 37461 13271 37519 13277
rect 37921 13311 37979 13317
rect 37921 13277 37933 13311
rect 37967 13277 37979 13311
rect 40494 13308 40500 13320
rect 40455 13280 40500 13308
rect 37921 13271 37979 13277
rect 37476 13240 37504 13271
rect 40494 13268 40500 13280
rect 40552 13268 40558 13320
rect 41138 13268 41144 13320
rect 41196 13308 41202 13320
rect 41233 13311 41291 13317
rect 41233 13308 41245 13311
rect 41196 13280 41245 13308
rect 41196 13268 41202 13280
rect 41233 13277 41245 13280
rect 41279 13277 41291 13311
rect 41233 13271 41291 13277
rect 41690 13268 41696 13320
rect 41748 13308 41754 13320
rect 41877 13311 41935 13317
rect 41877 13308 41889 13311
rect 41748 13280 41889 13308
rect 41748 13268 41754 13280
rect 41877 13277 41889 13280
rect 41923 13277 41935 13311
rect 41877 13271 41935 13277
rect 42794 13268 42800 13320
rect 42852 13308 42858 13320
rect 42889 13311 42947 13317
rect 42889 13308 42901 13311
rect 42852 13280 42901 13308
rect 42852 13268 42858 13280
rect 42889 13277 42901 13280
rect 42935 13277 42947 13311
rect 43530 13308 43536 13320
rect 43491 13280 43536 13308
rect 42889 13271 42947 13277
rect 43530 13268 43536 13280
rect 43588 13268 43594 13320
rect 41322 13240 41328 13252
rect 37476 13212 41328 13240
rect 41322 13200 41328 13212
rect 41380 13200 41386 13252
rect 42150 13240 42156 13252
rect 42063 13212 42156 13240
rect 42150 13200 42156 13212
rect 42208 13240 42214 13252
rect 43824 13240 43852 13475
rect 43990 13472 43996 13484
rect 44048 13472 44054 13524
rect 45462 13512 45468 13524
rect 44376 13484 45468 13512
rect 44269 13311 44327 13317
rect 44269 13277 44281 13311
rect 44315 13308 44327 13311
rect 44376 13308 44404 13484
rect 45462 13472 45468 13484
rect 45520 13512 45526 13524
rect 46109 13515 46167 13521
rect 46109 13512 46121 13515
rect 45520 13484 46121 13512
rect 45520 13472 45526 13484
rect 46109 13481 46121 13484
rect 46155 13481 46167 13515
rect 46109 13475 46167 13481
rect 52914 13472 52920 13524
rect 52972 13512 52978 13524
rect 53377 13515 53435 13521
rect 53377 13512 53389 13515
rect 52972 13484 53389 13512
rect 52972 13472 52978 13484
rect 53377 13481 53389 13484
rect 53423 13481 53435 13515
rect 53377 13475 53435 13481
rect 57974 13472 57980 13524
rect 58032 13512 58038 13524
rect 58161 13515 58219 13521
rect 58161 13512 58173 13515
rect 58032 13484 58173 13512
rect 58032 13472 58038 13484
rect 58161 13481 58173 13484
rect 58207 13481 58219 13515
rect 58161 13475 58219 13481
rect 49145 13447 49203 13453
rect 44468 13416 47348 13444
rect 44468 13317 44496 13416
rect 45186 13336 45192 13388
rect 45244 13376 45250 13388
rect 45281 13379 45339 13385
rect 45281 13376 45293 13379
rect 45244 13348 45293 13376
rect 45244 13336 45250 13348
rect 45281 13345 45293 13348
rect 45327 13345 45339 13379
rect 45281 13339 45339 13345
rect 45373 13379 45431 13385
rect 45373 13345 45385 13379
rect 45419 13376 45431 13379
rect 45419 13348 46336 13376
rect 45419 13345 45431 13348
rect 45373 13339 45431 13345
rect 46308 13320 46336 13348
rect 44315 13280 44404 13308
rect 44453 13311 44511 13317
rect 44315 13277 44327 13280
rect 44269 13271 44327 13277
rect 44453 13277 44465 13311
rect 44499 13277 44511 13311
rect 44453 13271 44511 13277
rect 44818 13268 44824 13320
rect 44876 13308 44882 13320
rect 45465 13311 45523 13317
rect 45465 13308 45477 13311
rect 44876 13280 45477 13308
rect 44876 13268 44882 13280
rect 45465 13277 45477 13280
rect 45511 13277 45523 13311
rect 45465 13271 45523 13277
rect 42208 13212 43852 13240
rect 44361 13243 44419 13249
rect 42208 13200 42214 13212
rect 44361 13209 44373 13243
rect 44407 13240 44419 13243
rect 45370 13240 45376 13252
rect 44407 13212 45376 13240
rect 44407 13209 44419 13212
rect 44361 13203 44419 13209
rect 45370 13200 45376 13212
rect 45428 13200 45434 13252
rect 45480 13240 45508 13271
rect 45554 13268 45560 13320
rect 45612 13308 45618 13320
rect 46290 13308 46296 13320
rect 45612 13280 45657 13308
rect 46251 13280 46296 13308
rect 45612 13268 45618 13280
rect 46290 13268 46296 13280
rect 46348 13268 46354 13320
rect 47210 13308 47216 13320
rect 47171 13280 47216 13308
rect 47210 13268 47216 13280
rect 47268 13268 47274 13320
rect 47320 13240 47348 13416
rect 49145 13413 49157 13447
rect 49191 13444 49203 13447
rect 50614 13444 50620 13456
rect 49191 13416 50620 13444
rect 49191 13413 49203 13416
rect 49145 13407 49203 13413
rect 50614 13404 50620 13416
rect 50672 13404 50678 13456
rect 50249 13379 50307 13385
rect 50249 13376 50261 13379
rect 47412 13348 50261 13376
rect 47412 13317 47440 13348
rect 50249 13345 50261 13348
rect 50295 13345 50307 13379
rect 51902 13376 51908 13388
rect 51863 13348 51908 13376
rect 50249 13339 50307 13345
rect 51902 13336 51908 13348
rect 51960 13336 51966 13388
rect 53374 13336 53380 13388
rect 53432 13376 53438 13388
rect 54205 13379 54263 13385
rect 54205 13376 54217 13379
rect 53432 13348 54217 13376
rect 53432 13336 53438 13348
rect 54205 13345 54217 13348
rect 54251 13345 54263 13379
rect 56686 13376 56692 13388
rect 56647 13348 56692 13376
rect 54205 13339 54263 13345
rect 56686 13336 56692 13348
rect 56744 13336 56750 13388
rect 47397 13311 47455 13317
rect 47397 13277 47409 13311
rect 47443 13277 47455 13311
rect 47397 13271 47455 13277
rect 47486 13268 47492 13320
rect 47544 13308 47550 13320
rect 48222 13308 48228 13320
rect 47544 13280 47637 13308
rect 48135 13280 48228 13308
rect 47544 13268 47550 13280
rect 48222 13268 48228 13280
rect 48280 13308 48286 13320
rect 50157 13311 50215 13317
rect 50157 13308 50169 13311
rect 48280 13280 50169 13308
rect 48280 13268 48286 13280
rect 50157 13277 50169 13280
rect 50203 13277 50215 13311
rect 50338 13308 50344 13320
rect 50299 13280 50344 13308
rect 50157 13271 50215 13277
rect 50338 13268 50344 13280
rect 50396 13268 50402 13320
rect 50798 13308 50804 13320
rect 50759 13280 50804 13308
rect 50798 13268 50804 13280
rect 50856 13268 50862 13320
rect 51350 13308 51356 13320
rect 51046 13280 51356 13308
rect 47504 13240 47532 13268
rect 48774 13240 48780 13252
rect 45480 13212 47164 13240
rect 47320 13212 47532 13240
rect 48735 13212 48780 13240
rect 34848 13144 37412 13172
rect 38105 13175 38163 13181
rect 34848 13132 34854 13144
rect 38105 13141 38117 13175
rect 38151 13172 38163 13175
rect 38194 13172 38200 13184
rect 38151 13144 38200 13172
rect 38151 13141 38163 13144
rect 38105 13135 38163 13141
rect 38194 13132 38200 13144
rect 38252 13132 38258 13184
rect 44910 13132 44916 13184
rect 44968 13172 44974 13184
rect 45097 13175 45155 13181
rect 45097 13172 45109 13175
rect 44968 13144 45109 13172
rect 44968 13132 44974 13144
rect 45097 13141 45109 13144
rect 45143 13141 45155 13175
rect 47026 13172 47032 13184
rect 46987 13144 47032 13172
rect 45097 13135 45155 13141
rect 47026 13132 47032 13144
rect 47084 13132 47090 13184
rect 47136 13172 47164 13212
rect 48774 13200 48780 13212
rect 48832 13200 48838 13252
rect 49786 13200 49792 13252
rect 49844 13240 49850 13252
rect 51046 13240 51074 13280
rect 51350 13268 51356 13280
rect 51408 13308 51414 13320
rect 51629 13311 51687 13317
rect 51629 13308 51641 13311
rect 51408 13280 51641 13308
rect 51408 13268 51414 13280
rect 51629 13277 51641 13280
rect 51675 13277 51687 13311
rect 51629 13271 51687 13277
rect 53558 13268 53564 13320
rect 53616 13308 53622 13320
rect 54297 13311 54355 13317
rect 54297 13308 54309 13311
rect 53616 13280 54309 13308
rect 53616 13268 53622 13280
rect 54297 13277 54309 13280
rect 54343 13277 54355 13311
rect 54297 13271 54355 13277
rect 55582 13268 55588 13320
rect 55640 13308 55646 13320
rect 56413 13311 56471 13317
rect 56413 13308 56425 13311
rect 55640 13280 56425 13308
rect 55640 13268 55646 13280
rect 56413 13277 56425 13280
rect 56459 13277 56471 13311
rect 56413 13271 56471 13277
rect 53190 13240 53196 13252
rect 49844 13212 51074 13240
rect 53130 13212 53196 13240
rect 49844 13200 49850 13212
rect 48133 13175 48191 13181
rect 48133 13172 48145 13175
rect 47136 13144 48145 13172
rect 48133 13141 48145 13144
rect 48179 13172 48191 13175
rect 48314 13172 48320 13184
rect 48179 13144 48320 13172
rect 48179 13141 48191 13144
rect 48133 13135 48191 13141
rect 48314 13132 48320 13144
rect 48372 13132 48378 13184
rect 49237 13175 49295 13181
rect 49237 13141 49249 13175
rect 49283 13172 49295 13175
rect 49326 13172 49332 13184
rect 49283 13144 49332 13172
rect 49283 13141 49295 13144
rect 49237 13135 49295 13141
rect 49326 13132 49332 13144
rect 49384 13132 49390 13184
rect 51000 13181 51028 13212
rect 53190 13200 53196 13212
rect 53248 13200 53254 13252
rect 57330 13200 57336 13252
rect 57388 13200 57394 13252
rect 50985 13175 51043 13181
rect 50985 13141 50997 13175
rect 51031 13172 51043 13175
rect 54665 13175 54723 13181
rect 51031 13144 51065 13172
rect 51031 13141 51043 13144
rect 50985 13135 51043 13141
rect 54665 13141 54677 13175
rect 54711 13172 54723 13175
rect 55306 13172 55312 13184
rect 54711 13144 55312 13172
rect 54711 13141 54723 13144
rect 54665 13135 54723 13141
rect 55306 13132 55312 13144
rect 55364 13132 55370 13184
rect 1104 13082 58880 13104
rect 1104 13030 15398 13082
rect 15450 13030 15462 13082
rect 15514 13030 15526 13082
rect 15578 13030 15590 13082
rect 15642 13030 15654 13082
rect 15706 13030 29846 13082
rect 29898 13030 29910 13082
rect 29962 13030 29974 13082
rect 30026 13030 30038 13082
rect 30090 13030 30102 13082
rect 30154 13030 44294 13082
rect 44346 13030 44358 13082
rect 44410 13030 44422 13082
rect 44474 13030 44486 13082
rect 44538 13030 44550 13082
rect 44602 13030 58880 13082
rect 1104 13008 58880 13030
rect 9674 12968 9680 12980
rect 9635 12940 9680 12968
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 16942 12968 16948 12980
rect 10100 12940 16948 12968
rect 10100 12928 10106 12940
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18322 12968 18328 12980
rect 18012 12940 18328 12968
rect 18012 12928 18018 12940
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 20901 12971 20959 12977
rect 20901 12937 20913 12971
rect 20947 12968 20959 12971
rect 22462 12968 22468 12980
rect 20947 12940 22468 12968
rect 20947 12937 20959 12940
rect 20901 12931 20959 12937
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 23198 12928 23204 12980
rect 23256 12968 23262 12980
rect 25777 12971 25835 12977
rect 25777 12968 25789 12971
rect 23256 12940 25789 12968
rect 23256 12928 23262 12940
rect 25777 12937 25789 12940
rect 25823 12937 25835 12971
rect 25777 12931 25835 12937
rect 26510 12928 26516 12980
rect 26568 12968 26574 12980
rect 26973 12971 27031 12977
rect 26973 12968 26985 12971
rect 26568 12940 26985 12968
rect 26568 12928 26574 12940
rect 26973 12937 26985 12940
rect 27019 12937 27031 12971
rect 26973 12931 27031 12937
rect 30282 12928 30288 12980
rect 30340 12968 30346 12980
rect 30837 12971 30895 12977
rect 30837 12968 30849 12971
rect 30340 12940 30849 12968
rect 30340 12928 30346 12940
rect 30837 12937 30849 12940
rect 30883 12937 30895 12971
rect 30837 12931 30895 12937
rect 31005 12971 31063 12977
rect 31005 12937 31017 12971
rect 31051 12968 31063 12971
rect 31110 12968 31116 12980
rect 31051 12940 31116 12968
rect 31051 12937 31063 12940
rect 31005 12931 31063 12937
rect 31110 12928 31116 12940
rect 31168 12928 31174 12980
rect 35342 12968 35348 12980
rect 33520 12940 35348 12968
rect 10962 12900 10968 12912
rect 10923 12872 10968 12900
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 14366 12900 14372 12912
rect 14327 12872 14372 12900
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 17310 12900 17316 12912
rect 17271 12872 17316 12900
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 19978 12860 19984 12912
rect 20036 12900 20042 12912
rect 22373 12903 22431 12909
rect 22373 12900 22385 12903
rect 20036 12872 22385 12900
rect 20036 12860 20042 12872
rect 22373 12869 22385 12872
rect 22419 12869 22431 12903
rect 23750 12900 23756 12912
rect 23598 12872 23756 12900
rect 22373 12863 22431 12869
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 24210 12860 24216 12912
rect 24268 12900 24274 12912
rect 24489 12903 24547 12909
rect 24489 12900 24501 12903
rect 24268 12872 24501 12900
rect 24268 12860 24274 12872
rect 24489 12869 24501 12872
rect 24535 12869 24547 12903
rect 29454 12900 29460 12912
rect 24489 12863 24547 12869
rect 27724 12872 29460 12900
rect 7466 12792 7472 12844
rect 7524 12832 7530 12844
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 7524 12804 7665 12832
rect 7524 12792 7530 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11204 12804 11805 12832
rect 11204 12792 11210 12804
rect 11793 12801 11805 12804
rect 11839 12832 11851 12835
rect 11882 12832 11888 12844
rect 11839 12804 11888 12832
rect 11839 12801 11851 12804
rect 11793 12795 11851 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 12066 12832 12072 12844
rect 12027 12804 12072 12832
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12618 12832 12624 12844
rect 12579 12804 12624 12832
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 13538 12832 13544 12844
rect 13499 12804 13544 12832
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 19886 12832 19892 12844
rect 19847 12804 19892 12832
rect 19886 12792 19892 12804
rect 19944 12792 19950 12844
rect 20257 12835 20315 12841
rect 20257 12801 20269 12835
rect 20303 12832 20315 12835
rect 22094 12832 22100 12844
rect 20303 12804 21128 12832
rect 22055 12804 22100 12832
rect 20303 12801 20315 12804
rect 20257 12795 20315 12801
rect 7742 12764 7748 12776
rect 7703 12736 7748 12764
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13504 12736 13645 12764
rect 13504 12724 13510 12736
rect 13633 12733 13645 12736
rect 13679 12764 13691 12767
rect 13722 12764 13728 12776
rect 13679 12736 13728 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 17034 12764 17040 12776
rect 16163 12736 17040 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12733 17187 12767
rect 18598 12764 18604 12776
rect 18559 12736 18604 12764
rect 17129 12727 17187 12733
rect 13909 12699 13967 12705
rect 13909 12665 13921 12699
rect 13955 12696 13967 12699
rect 15010 12696 15016 12708
rect 13955 12668 15016 12696
rect 13955 12665 13967 12668
rect 13909 12659 13967 12665
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 17144 12696 17172 12727
rect 18598 12724 18604 12736
rect 18656 12764 18662 12776
rect 18966 12764 18972 12776
rect 18656 12736 18972 12764
rect 18656 12724 18662 12736
rect 18966 12724 18972 12736
rect 19024 12724 19030 12776
rect 21100 12764 21128 12804
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 27724 12841 27752 12872
rect 29454 12860 29460 12872
rect 29512 12860 29518 12912
rect 29822 12900 29828 12912
rect 29783 12872 29828 12900
rect 29822 12860 29828 12872
rect 29880 12860 29886 12912
rect 31202 12900 31208 12912
rect 31163 12872 31208 12900
rect 31202 12860 31208 12872
rect 31260 12860 31266 12912
rect 27709 12835 27767 12841
rect 27709 12801 27721 12835
rect 27755 12801 27767 12835
rect 27709 12795 27767 12801
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12832 32367 12835
rect 33520 12832 33548 12940
rect 35342 12928 35348 12940
rect 35400 12928 35406 12980
rect 35526 12968 35532 12980
rect 35487 12940 35532 12968
rect 35526 12928 35532 12940
rect 35584 12928 35590 12980
rect 39390 12928 39396 12980
rect 39448 12968 39454 12980
rect 40954 12968 40960 12980
rect 39448 12940 40960 12968
rect 39448 12928 39454 12940
rect 40954 12928 40960 12940
rect 41012 12928 41018 12980
rect 41690 12928 41696 12980
rect 41748 12968 41754 12980
rect 42613 12971 42671 12977
rect 42613 12968 42625 12971
rect 41748 12940 42625 12968
rect 41748 12928 41754 12940
rect 42613 12937 42625 12940
rect 42659 12937 42671 12971
rect 48774 12968 48780 12980
rect 42613 12931 42671 12937
rect 45112 12940 48780 12968
rect 34790 12860 34796 12912
rect 34848 12860 34854 12912
rect 45112 12900 45140 12940
rect 48774 12928 48780 12940
rect 48832 12968 48838 12980
rect 50341 12971 50399 12977
rect 50341 12968 50353 12971
rect 48832 12940 50353 12968
rect 48832 12928 48838 12940
rect 50341 12937 50353 12940
rect 50387 12968 50399 12971
rect 50430 12968 50436 12980
rect 50387 12940 50436 12968
rect 50387 12937 50399 12940
rect 50341 12931 50399 12937
rect 50430 12928 50436 12940
rect 50488 12928 50494 12980
rect 53190 12968 53196 12980
rect 50540 12940 53196 12968
rect 37292 12872 45140 12900
rect 45572 12872 49464 12900
rect 32355 12804 33548 12832
rect 32355 12801 32367 12804
rect 32309 12795 32367 12801
rect 33594 12792 33600 12844
rect 33652 12832 33658 12844
rect 33778 12832 33784 12844
rect 33652 12804 33784 12832
rect 33652 12792 33658 12804
rect 33778 12792 33784 12804
rect 33836 12792 33842 12844
rect 35986 12832 35992 12844
rect 35947 12804 35992 12832
rect 35986 12792 35992 12804
rect 36044 12792 36050 12844
rect 37292 12841 37320 12872
rect 37277 12835 37335 12841
rect 37277 12801 37289 12835
rect 37323 12801 37335 12835
rect 37277 12795 37335 12801
rect 39117 12835 39175 12841
rect 39117 12801 39129 12835
rect 39163 12832 39175 12835
rect 39390 12832 39396 12844
rect 39163 12804 39396 12832
rect 39163 12801 39175 12804
rect 39117 12795 39175 12801
rect 39390 12792 39396 12804
rect 39448 12792 39454 12844
rect 40586 12792 40592 12844
rect 40644 12832 40650 12844
rect 40681 12835 40739 12841
rect 40681 12832 40693 12835
rect 40644 12804 40693 12832
rect 40644 12792 40650 12804
rect 40681 12801 40693 12804
rect 40727 12801 40739 12835
rect 40954 12832 40960 12844
rect 40915 12804 40960 12832
rect 40681 12795 40739 12801
rect 40954 12792 40960 12804
rect 41012 12792 41018 12844
rect 41693 12835 41751 12841
rect 41693 12801 41705 12835
rect 41739 12832 41751 12835
rect 42429 12835 42487 12841
rect 42429 12832 42441 12835
rect 41739 12804 42441 12832
rect 41739 12801 41751 12804
rect 41693 12795 41751 12801
rect 42429 12801 42441 12804
rect 42475 12832 42487 12835
rect 43530 12832 43536 12844
rect 42475 12804 43536 12832
rect 42475 12801 42487 12804
rect 42429 12795 42487 12801
rect 43530 12792 43536 12804
rect 43588 12792 43594 12844
rect 44269 12835 44327 12841
rect 44269 12801 44281 12835
rect 44315 12832 44327 12835
rect 44726 12832 44732 12844
rect 44315 12804 44732 12832
rect 44315 12801 44327 12804
rect 44269 12795 44327 12801
rect 44726 12792 44732 12804
rect 44784 12792 44790 12844
rect 44910 12832 44916 12844
rect 44871 12804 44916 12832
rect 44910 12792 44916 12804
rect 44968 12792 44974 12844
rect 45186 12792 45192 12844
rect 45244 12832 45250 12844
rect 45465 12835 45523 12841
rect 45465 12832 45477 12835
rect 45244 12804 45477 12832
rect 45244 12792 45250 12804
rect 45465 12801 45477 12804
rect 45511 12801 45523 12835
rect 45465 12795 45523 12801
rect 23014 12764 23020 12776
rect 21100 12736 23020 12764
rect 23014 12724 23020 12736
rect 23072 12724 23078 12776
rect 28169 12767 28227 12773
rect 28169 12764 28181 12767
rect 23400 12736 28181 12764
rect 18138 12696 18144 12708
rect 17144 12668 18144 12696
rect 18138 12656 18144 12668
rect 18196 12656 18202 12708
rect 18984 12696 19012 12724
rect 18984 12668 22094 12696
rect 7926 12628 7932 12640
rect 7887 12600 7932 12628
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 14274 12588 14280 12640
rect 14332 12628 14338 12640
rect 17126 12628 17132 12640
rect 14332 12600 17132 12628
rect 14332 12588 14338 12600
rect 17126 12588 17132 12600
rect 17184 12588 17190 12640
rect 22066 12628 22094 12668
rect 23400 12628 23428 12736
rect 28169 12733 28181 12736
rect 28215 12733 28227 12767
rect 28169 12727 28227 12733
rect 30009 12767 30067 12773
rect 30009 12733 30021 12767
rect 30055 12733 30067 12767
rect 32214 12764 32220 12776
rect 32175 12736 32220 12764
rect 30009 12727 30067 12733
rect 23842 12628 23848 12640
rect 22066 12600 23428 12628
rect 23803 12600 23848 12628
rect 23842 12588 23848 12600
rect 23900 12588 23906 12640
rect 27614 12628 27620 12640
rect 27575 12600 27620 12628
rect 27614 12588 27620 12600
rect 27672 12588 27678 12640
rect 28184 12628 28212 12727
rect 30024 12696 30052 12727
rect 32214 12724 32220 12736
rect 32272 12724 32278 12776
rect 33134 12764 33140 12776
rect 33095 12736 33140 12764
rect 33134 12724 33140 12736
rect 33192 12724 33198 12776
rect 34054 12764 34060 12776
rect 34015 12736 34060 12764
rect 34054 12724 34060 12736
rect 34112 12724 34118 12776
rect 35526 12724 35532 12776
rect 35584 12764 35590 12776
rect 36081 12767 36139 12773
rect 36081 12764 36093 12767
rect 35584 12736 36093 12764
rect 35584 12724 35590 12736
rect 36081 12733 36093 12736
rect 36127 12733 36139 12767
rect 37458 12764 37464 12776
rect 37419 12736 37464 12764
rect 36081 12727 36139 12733
rect 37458 12724 37464 12736
rect 37516 12724 37522 12776
rect 40126 12764 40132 12776
rect 40087 12736 40132 12764
rect 40126 12724 40132 12736
rect 40184 12724 40190 12776
rect 41877 12767 41935 12773
rect 41877 12733 41889 12767
rect 41923 12764 41935 12767
rect 42150 12764 42156 12776
rect 41923 12736 42156 12764
rect 41923 12733 41935 12736
rect 41877 12727 41935 12733
rect 42150 12724 42156 12736
rect 42208 12724 42214 12776
rect 45278 12724 45284 12776
rect 45336 12764 45342 12776
rect 45572 12764 45600 12872
rect 46750 12792 46756 12844
rect 46808 12832 46814 12844
rect 46845 12835 46903 12841
rect 46845 12832 46857 12835
rect 46808 12804 46857 12832
rect 46808 12792 46814 12804
rect 46845 12801 46857 12804
rect 46891 12801 46903 12835
rect 46845 12795 46903 12801
rect 48222 12792 48228 12844
rect 48280 12832 48286 12844
rect 48317 12835 48375 12841
rect 48317 12832 48329 12835
rect 48280 12804 48329 12832
rect 48280 12792 48286 12804
rect 48317 12801 48329 12804
rect 48363 12801 48375 12835
rect 49326 12832 49332 12844
rect 49287 12804 49332 12832
rect 48317 12795 48375 12801
rect 49326 12792 49332 12804
rect 49384 12792 49390 12844
rect 49436 12841 49464 12872
rect 50246 12860 50252 12912
rect 50304 12900 50310 12912
rect 50540 12900 50568 12940
rect 53190 12928 53196 12940
rect 53248 12928 53254 12980
rect 53374 12968 53380 12980
rect 53335 12940 53380 12968
rect 53374 12928 53380 12940
rect 53432 12928 53438 12980
rect 53558 12928 53564 12980
rect 53616 12968 53622 12980
rect 53837 12971 53895 12977
rect 53837 12968 53849 12971
rect 53616 12940 53849 12968
rect 53616 12928 53622 12940
rect 53837 12937 53849 12940
rect 53883 12937 53895 12971
rect 55674 12968 55680 12980
rect 53837 12931 53895 12937
rect 54956 12940 55680 12968
rect 51813 12903 51871 12909
rect 50304 12872 50646 12900
rect 50304 12860 50310 12872
rect 51813 12869 51825 12903
rect 51859 12900 51871 12903
rect 51902 12900 51908 12912
rect 51859 12872 51908 12900
rect 51859 12869 51871 12872
rect 51813 12863 51871 12869
rect 51902 12860 51908 12872
rect 51960 12860 51966 12912
rect 54956 12900 54984 12940
rect 55674 12928 55680 12940
rect 55732 12928 55738 12980
rect 57333 12971 57391 12977
rect 57333 12937 57345 12971
rect 57379 12937 57391 12971
rect 58066 12968 58072 12980
rect 58027 12940 58072 12968
rect 57333 12931 57391 12937
rect 55306 12900 55312 12912
rect 54878 12872 54984 12900
rect 55267 12872 55312 12900
rect 55306 12860 55312 12872
rect 55364 12860 55370 12912
rect 55600 12872 57192 12900
rect 55600 12844 55628 12872
rect 57164 12844 57192 12872
rect 49421 12835 49479 12841
rect 49421 12801 49433 12835
rect 49467 12832 49479 12835
rect 50338 12832 50344 12844
rect 49467 12804 50344 12832
rect 49467 12801 49479 12804
rect 49421 12795 49479 12801
rect 50338 12792 50344 12804
rect 50396 12792 50402 12844
rect 53006 12792 53012 12844
rect 53064 12832 53070 12844
rect 53101 12835 53159 12841
rect 53101 12832 53113 12835
rect 53064 12804 53113 12832
rect 53064 12792 53070 12804
rect 53101 12801 53113 12804
rect 53147 12801 53159 12835
rect 53101 12795 53159 12801
rect 55582 12792 55588 12844
rect 55640 12832 55646 12844
rect 55640 12804 55685 12832
rect 55640 12792 55646 12804
rect 56042 12792 56048 12844
rect 56100 12832 56106 12844
rect 56137 12835 56195 12841
rect 56137 12832 56149 12835
rect 56100 12804 56149 12832
rect 56100 12792 56106 12804
rect 56137 12801 56149 12804
rect 56183 12801 56195 12835
rect 57146 12832 57152 12844
rect 57059 12804 57152 12832
rect 56137 12795 56195 12801
rect 57146 12792 57152 12804
rect 57204 12792 57210 12844
rect 57348 12832 57376 12931
rect 58066 12928 58072 12940
rect 58124 12928 58130 12980
rect 57885 12835 57943 12841
rect 57885 12832 57897 12835
rect 57348 12804 57897 12832
rect 57885 12801 57897 12804
rect 57931 12801 57943 12835
rect 57885 12795 57943 12801
rect 45336 12736 45600 12764
rect 45649 12767 45707 12773
rect 45336 12724 45342 12736
rect 45649 12733 45661 12767
rect 45695 12764 45707 12767
rect 48130 12764 48136 12776
rect 45695 12736 48136 12764
rect 45695 12733 45707 12736
rect 45649 12727 45707 12733
rect 48130 12724 48136 12736
rect 48188 12724 48194 12776
rect 48409 12767 48467 12773
rect 48409 12733 48421 12767
rect 48455 12764 48467 12767
rect 49142 12764 49148 12776
rect 48455 12736 48820 12764
rect 49103 12736 49148 12764
rect 48455 12733 48467 12736
rect 48409 12727 48467 12733
rect 32677 12699 32735 12705
rect 30024 12668 32628 12696
rect 30926 12628 30932 12640
rect 28184 12600 30932 12628
rect 30926 12588 30932 12600
rect 30984 12588 30990 12640
rect 31021 12631 31079 12637
rect 31021 12597 31033 12631
rect 31067 12628 31079 12631
rect 31478 12628 31484 12640
rect 31067 12600 31484 12628
rect 31067 12597 31079 12600
rect 31021 12591 31079 12597
rect 31478 12588 31484 12600
rect 31536 12628 31542 12640
rect 31662 12628 31668 12640
rect 31536 12600 31668 12628
rect 31536 12588 31542 12600
rect 31662 12588 31668 12600
rect 31720 12588 31726 12640
rect 32600 12628 32628 12668
rect 32677 12665 32689 12699
rect 32723 12696 32735 12699
rect 33226 12696 33232 12708
rect 32723 12668 33232 12696
rect 32723 12665 32735 12668
rect 32677 12659 32735 12665
rect 33226 12656 33232 12668
rect 33284 12656 33290 12708
rect 37642 12696 37648 12708
rect 35084 12668 37648 12696
rect 35084 12628 35112 12668
rect 37642 12656 37648 12668
rect 37700 12656 37706 12708
rect 41506 12656 41512 12708
rect 41564 12696 41570 12708
rect 46385 12699 46443 12705
rect 46385 12696 46397 12699
rect 41564 12668 46397 12696
rect 41564 12656 41570 12668
rect 46385 12665 46397 12668
rect 46431 12696 46443 12699
rect 46934 12696 46940 12708
rect 46431 12668 46940 12696
rect 46431 12665 46443 12668
rect 46385 12659 46443 12665
rect 46934 12656 46940 12668
rect 46992 12656 46998 12708
rect 47029 12699 47087 12705
rect 47029 12665 47041 12699
rect 47075 12696 47087 12699
rect 48682 12696 48688 12708
rect 47075 12668 48452 12696
rect 48643 12668 48688 12696
rect 47075 12665 47087 12668
rect 47029 12659 47087 12665
rect 48424 12640 48452 12668
rect 48682 12656 48688 12668
rect 48740 12656 48746 12708
rect 48792 12696 48820 12736
rect 49142 12724 49148 12736
rect 49200 12764 49206 12776
rect 49200 12736 50476 12764
rect 49200 12724 49206 12736
rect 49237 12699 49295 12705
rect 49237 12696 49249 12699
rect 48792 12668 49249 12696
rect 49237 12665 49249 12668
rect 49283 12665 49295 12699
rect 49237 12659 49295 12665
rect 32600 12600 35112 12628
rect 35434 12588 35440 12640
rect 35492 12628 35498 12640
rect 35989 12631 36047 12637
rect 35989 12628 36001 12631
rect 35492 12600 36001 12628
rect 35492 12588 35498 12600
rect 35989 12597 36001 12600
rect 36035 12597 36047 12631
rect 35989 12591 36047 12597
rect 36357 12631 36415 12637
rect 36357 12597 36369 12631
rect 36403 12628 36415 12631
rect 38470 12628 38476 12640
rect 36403 12600 38476 12628
rect 36403 12597 36415 12600
rect 36357 12591 36415 12597
rect 38470 12588 38476 12600
rect 38528 12588 38534 12640
rect 39669 12631 39727 12637
rect 39669 12597 39681 12631
rect 39715 12628 39727 12631
rect 40126 12628 40132 12640
rect 39715 12600 40132 12628
rect 39715 12597 39727 12600
rect 39669 12591 39727 12597
rect 40126 12588 40132 12600
rect 40184 12588 40190 12640
rect 44821 12631 44879 12637
rect 44821 12597 44833 12631
rect 44867 12628 44879 12631
rect 45278 12628 45284 12640
rect 44867 12600 45284 12628
rect 44867 12597 44879 12600
rect 44821 12591 44879 12597
rect 45278 12588 45284 12600
rect 45336 12588 45342 12640
rect 46474 12588 46480 12640
rect 46532 12628 46538 12640
rect 47581 12631 47639 12637
rect 47581 12628 47593 12631
rect 46532 12600 47593 12628
rect 46532 12588 46538 12600
rect 47581 12597 47593 12600
rect 47627 12597 47639 12631
rect 47581 12591 47639 12597
rect 48406 12588 48412 12640
rect 48464 12588 48470 12640
rect 50448 12628 50476 12736
rect 50798 12724 50804 12776
rect 50856 12764 50862 12776
rect 52089 12767 52147 12773
rect 52089 12764 52101 12767
rect 50856 12736 52101 12764
rect 50856 12724 50862 12736
rect 52089 12733 52101 12736
rect 52135 12733 52147 12767
rect 53374 12764 53380 12776
rect 53335 12736 53380 12764
rect 52089 12727 52147 12733
rect 53374 12724 53380 12736
rect 53432 12724 53438 12776
rect 55674 12724 55680 12776
rect 55732 12764 55738 12776
rect 56060 12764 56088 12792
rect 55732 12736 56088 12764
rect 55732 12724 55738 12736
rect 53193 12699 53251 12705
rect 53193 12665 53205 12699
rect 53239 12696 53251 12699
rect 53926 12696 53932 12708
rect 53239 12668 53932 12696
rect 53239 12665 53251 12668
rect 53193 12659 53251 12665
rect 53926 12656 53932 12668
rect 53984 12656 53990 12708
rect 56321 12699 56379 12705
rect 56321 12665 56333 12699
rect 56367 12696 56379 12699
rect 56594 12696 56600 12708
rect 56367 12668 56600 12696
rect 56367 12665 56379 12668
rect 56321 12659 56379 12665
rect 56594 12656 56600 12668
rect 56652 12656 56658 12708
rect 52362 12628 52368 12640
rect 50448 12600 52368 12628
rect 52362 12588 52368 12600
rect 52420 12588 52426 12640
rect 1104 12538 58880 12560
rect 1104 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 8302 12538
rect 8354 12486 8366 12538
rect 8418 12486 8430 12538
rect 8482 12486 22622 12538
rect 22674 12486 22686 12538
rect 22738 12486 22750 12538
rect 22802 12486 22814 12538
rect 22866 12486 22878 12538
rect 22930 12486 37070 12538
rect 37122 12486 37134 12538
rect 37186 12486 37198 12538
rect 37250 12486 37262 12538
rect 37314 12486 37326 12538
rect 37378 12486 51518 12538
rect 51570 12486 51582 12538
rect 51634 12486 51646 12538
rect 51698 12486 51710 12538
rect 51762 12486 51774 12538
rect 51826 12486 58880 12538
rect 1104 12464 58880 12486
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 10873 12427 10931 12433
rect 10873 12424 10885 12427
rect 10836 12396 10885 12424
rect 10836 12384 10842 12396
rect 10873 12393 10885 12396
rect 10919 12393 10931 12427
rect 10873 12387 10931 12393
rect 14185 12427 14243 12433
rect 14185 12393 14197 12427
rect 14231 12424 14243 12427
rect 14734 12424 14740 12436
rect 14231 12396 14740 12424
rect 14231 12393 14243 12396
rect 14185 12387 14243 12393
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 15105 12427 15163 12433
rect 15105 12393 15117 12427
rect 15151 12424 15163 12427
rect 16758 12424 16764 12436
rect 15151 12396 16764 12424
rect 15151 12393 15163 12396
rect 15105 12387 15163 12393
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 16850 12384 16856 12436
rect 16908 12424 16914 12436
rect 19426 12424 19432 12436
rect 16908 12396 19432 12424
rect 16908 12384 16914 12396
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 23750 12424 23756 12436
rect 23711 12396 23756 12424
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 24397 12427 24455 12433
rect 24397 12393 24409 12427
rect 24443 12393 24455 12427
rect 24397 12387 24455 12393
rect 18230 12356 18236 12368
rect 16868 12328 18236 12356
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13354 12288 13360 12300
rect 13311 12260 13360 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 12676 12192 13185 12220
rect 12676 12180 12682 12192
rect 13173 12189 13185 12192
rect 13219 12220 13231 12223
rect 13538 12220 13544 12232
rect 13219 12192 13544 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 16868 12229 16896 12328
rect 18230 12316 18236 12328
rect 18288 12316 18294 12368
rect 18322 12316 18328 12368
rect 18380 12356 18386 12368
rect 18380 12328 19472 12356
rect 18380 12316 18386 12328
rect 19444 12288 19472 12328
rect 19518 12316 19524 12368
rect 19576 12356 19582 12368
rect 20254 12356 20260 12368
rect 19576 12328 20260 12356
rect 19576 12316 19582 12328
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 21269 12359 21327 12365
rect 21269 12325 21281 12359
rect 21315 12325 21327 12359
rect 21269 12319 21327 12325
rect 21284 12288 21312 12319
rect 21358 12316 21364 12368
rect 21416 12356 21422 12368
rect 24412 12356 24440 12387
rect 30374 12384 30380 12436
rect 30432 12424 30438 12436
rect 30469 12427 30527 12433
rect 30469 12424 30481 12427
rect 30432 12396 30481 12424
rect 30432 12384 30438 12396
rect 30469 12393 30481 12396
rect 30515 12393 30527 12427
rect 30469 12387 30527 12393
rect 30650 12384 30656 12436
rect 30708 12424 30714 12436
rect 31021 12427 31079 12433
rect 31021 12424 31033 12427
rect 30708 12396 31033 12424
rect 30708 12384 30714 12396
rect 31021 12393 31033 12396
rect 31067 12424 31079 12427
rect 31294 12424 31300 12436
rect 31067 12396 31300 12424
rect 31067 12393 31079 12396
rect 31021 12387 31079 12393
rect 31294 12384 31300 12396
rect 31352 12384 31358 12436
rect 31386 12384 31392 12436
rect 31444 12424 31450 12436
rect 33686 12424 33692 12436
rect 31444 12396 33692 12424
rect 31444 12384 31450 12396
rect 33686 12384 33692 12396
rect 33744 12384 33750 12436
rect 38746 12384 38752 12436
rect 38804 12424 38810 12436
rect 39301 12427 39359 12433
rect 39301 12424 39313 12427
rect 38804 12396 39313 12424
rect 38804 12384 38810 12396
rect 39301 12393 39313 12396
rect 39347 12424 39359 12427
rect 41506 12424 41512 12436
rect 39347 12396 41512 12424
rect 39347 12393 39359 12396
rect 39301 12387 39359 12393
rect 41506 12384 41512 12396
rect 41564 12384 41570 12436
rect 42150 12424 42156 12436
rect 42111 12396 42156 12424
rect 42150 12384 42156 12396
rect 42208 12384 42214 12436
rect 46290 12424 46296 12436
rect 43916 12396 46296 12424
rect 21416 12328 24440 12356
rect 28721 12359 28779 12365
rect 21416 12316 21422 12328
rect 28721 12325 28733 12359
rect 28767 12356 28779 12359
rect 29086 12356 29092 12368
rect 28767 12328 29092 12356
rect 28767 12325 28779 12328
rect 28721 12319 28779 12325
rect 29086 12316 29092 12328
rect 29144 12316 29150 12368
rect 30282 12356 30288 12368
rect 30243 12328 30288 12356
rect 30282 12316 30288 12328
rect 30340 12316 30346 12368
rect 31202 12316 31208 12368
rect 31260 12356 31266 12368
rect 34054 12356 34060 12368
rect 31260 12328 33916 12356
rect 34015 12328 34060 12356
rect 31260 12316 31266 12328
rect 24394 12288 24400 12300
rect 19444 12260 21220 12288
rect 21284 12260 24400 12288
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12220 18751 12223
rect 18966 12220 18972 12232
rect 18739 12192 18972 12220
rect 18739 12189 18751 12192
rect 18693 12183 18751 12189
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 19337 12223 19395 12229
rect 19337 12189 19349 12223
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 21082 12220 21088 12232
rect 19751 12192 21088 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 12161 12155 12219 12161
rect 12161 12121 12173 12155
rect 12207 12152 12219 12155
rect 13078 12152 13084 12164
rect 12207 12124 13084 12152
rect 12207 12121 12219 12124
rect 12161 12115 12219 12121
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 16390 12152 16396 12164
rect 16351 12124 16396 12152
rect 16390 12112 16396 12124
rect 16448 12112 16454 12164
rect 17037 12155 17095 12161
rect 17037 12121 17049 12155
rect 17083 12121 17095 12155
rect 17037 12115 17095 12121
rect 13538 12084 13544 12096
rect 13499 12056 13544 12084
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17052 12084 17080 12115
rect 17126 12112 17132 12164
rect 17184 12152 17190 12164
rect 19352 12152 19380 12183
rect 21082 12180 21088 12192
rect 21140 12180 21146 12232
rect 21192 12220 21220 12260
rect 21818 12220 21824 12232
rect 21192 12192 21824 12220
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 23860 12229 23888 12260
rect 24394 12248 24400 12260
rect 24452 12248 24458 12300
rect 24578 12248 24584 12300
rect 24636 12288 24642 12300
rect 25869 12291 25927 12297
rect 25869 12288 25881 12291
rect 24636 12260 25881 12288
rect 24636 12248 24642 12260
rect 25869 12257 25881 12260
rect 25915 12257 25927 12291
rect 25869 12251 25927 12257
rect 28445 12291 28503 12297
rect 28445 12257 28457 12291
rect 28491 12288 28503 12291
rect 28626 12288 28632 12300
rect 28491 12260 28632 12288
rect 28491 12257 28503 12260
rect 28445 12251 28503 12257
rect 28626 12248 28632 12260
rect 28684 12248 28690 12300
rect 29546 12248 29552 12300
rect 29604 12288 29610 12300
rect 32217 12291 32275 12297
rect 32217 12288 32229 12291
rect 29604 12260 32229 12288
rect 29604 12248 29610 12260
rect 32217 12257 32229 12260
rect 32263 12257 32275 12291
rect 32217 12251 32275 12257
rect 33410 12248 33416 12300
rect 33468 12288 33474 12300
rect 33597 12291 33655 12297
rect 33597 12288 33609 12291
rect 33468 12260 33609 12288
rect 33468 12248 33474 12260
rect 33597 12257 33609 12260
rect 33643 12257 33655 12291
rect 33597 12251 33655 12257
rect 23017 12223 23075 12229
rect 23017 12220 23029 12223
rect 21928 12192 23029 12220
rect 21928 12152 21956 12192
rect 23017 12189 23029 12192
rect 23063 12189 23075 12223
rect 23017 12183 23075 12189
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 26142 12180 26148 12232
rect 26200 12220 26206 12232
rect 26200 12192 26245 12220
rect 26200 12180 26206 12192
rect 26418 12180 26424 12232
rect 26476 12220 26482 12232
rect 26697 12223 26755 12229
rect 26697 12220 26709 12223
rect 26476 12192 26709 12220
rect 26476 12180 26482 12192
rect 26697 12189 26709 12192
rect 26743 12189 26755 12223
rect 26878 12220 26884 12232
rect 26839 12192 26884 12220
rect 26697 12183 26755 12189
rect 26878 12180 26884 12192
rect 26936 12180 26942 12232
rect 28353 12223 28411 12229
rect 28353 12189 28365 12223
rect 28399 12220 28411 12223
rect 30009 12223 30067 12229
rect 30009 12220 30021 12223
rect 28399 12192 30021 12220
rect 28399 12189 28411 12192
rect 28353 12183 28411 12189
rect 30009 12189 30021 12192
rect 30055 12220 30067 12223
rect 30650 12220 30656 12232
rect 30055 12192 30656 12220
rect 30055 12189 30067 12192
rect 30009 12183 30067 12189
rect 30650 12180 30656 12192
rect 30708 12180 30714 12232
rect 31202 12220 31208 12232
rect 31163 12192 31208 12220
rect 31202 12180 31208 12192
rect 31260 12180 31266 12232
rect 31297 12223 31355 12229
rect 31297 12189 31309 12223
rect 31343 12220 31355 12223
rect 31941 12223 31999 12229
rect 31941 12220 31953 12223
rect 31343 12192 31953 12220
rect 31343 12189 31355 12192
rect 31297 12183 31355 12189
rect 31941 12189 31953 12192
rect 31987 12189 31999 12223
rect 33686 12220 33692 12232
rect 33647 12192 33692 12220
rect 31941 12183 31999 12189
rect 17184 12124 21956 12152
rect 17184 12112 17190 12124
rect 22094 12112 22100 12164
rect 22152 12152 22158 12164
rect 22557 12155 22615 12161
rect 22557 12152 22569 12155
rect 22152 12124 22569 12152
rect 22152 12112 22158 12124
rect 22557 12121 22569 12124
rect 22603 12152 22615 12155
rect 23198 12152 23204 12164
rect 22603 12124 23204 12152
rect 22603 12121 22615 12124
rect 22557 12115 22615 12121
rect 23198 12112 23204 12124
rect 23256 12112 23262 12164
rect 25406 12112 25412 12164
rect 25464 12112 25470 12164
rect 31018 12152 31024 12164
rect 30979 12124 31024 12152
rect 31018 12112 31024 12124
rect 31076 12112 31082 12164
rect 31956 12152 31984 12183
rect 33686 12180 33692 12192
rect 33744 12180 33750 12232
rect 33888 12220 33916 12328
rect 34054 12316 34060 12328
rect 34112 12316 34118 12368
rect 36906 12316 36912 12368
rect 36964 12356 36970 12368
rect 37185 12359 37243 12365
rect 37185 12356 37197 12359
rect 36964 12328 37197 12356
rect 36964 12316 36970 12328
rect 37185 12325 37197 12328
rect 37231 12325 37243 12359
rect 39850 12356 39856 12368
rect 37185 12319 37243 12325
rect 38304 12328 39856 12356
rect 34790 12288 34796 12300
rect 34751 12260 34796 12288
rect 34790 12248 34796 12260
rect 34848 12248 34854 12300
rect 35437 12291 35495 12297
rect 35437 12257 35449 12291
rect 35483 12288 35495 12291
rect 35894 12288 35900 12300
rect 35483 12260 35900 12288
rect 35483 12257 35495 12260
rect 35437 12251 35495 12257
rect 35894 12248 35900 12260
rect 35952 12288 35958 12300
rect 36354 12288 36360 12300
rect 35952 12260 36360 12288
rect 35952 12248 35958 12260
rect 36354 12248 36360 12260
rect 36412 12248 36418 12300
rect 37645 12291 37703 12297
rect 37645 12257 37657 12291
rect 37691 12288 37703 12291
rect 38197 12291 38255 12297
rect 38197 12288 38209 12291
rect 37691 12260 38209 12288
rect 37691 12257 37703 12260
rect 37645 12251 37703 12257
rect 38197 12257 38209 12260
rect 38243 12257 38255 12291
rect 38197 12251 38255 12257
rect 34701 12223 34759 12229
rect 34701 12220 34713 12223
rect 33888 12192 34713 12220
rect 34701 12189 34713 12192
rect 34747 12189 34759 12223
rect 34882 12220 34888 12232
rect 34843 12192 34888 12220
rect 34701 12183 34759 12189
rect 34514 12152 34520 12164
rect 31956 12124 34520 12152
rect 34514 12112 34520 12124
rect 34572 12112 34578 12164
rect 34716 12152 34744 12183
rect 34882 12180 34888 12192
rect 34940 12180 34946 12232
rect 35713 12223 35771 12229
rect 35713 12189 35725 12223
rect 35759 12189 35771 12223
rect 35713 12183 35771 12189
rect 35728 12152 35756 12183
rect 36262 12180 36268 12232
rect 36320 12220 36326 12232
rect 37553 12223 37611 12229
rect 37553 12220 37565 12223
rect 36320 12192 37565 12220
rect 36320 12180 36326 12192
rect 37553 12189 37565 12192
rect 37599 12189 37611 12223
rect 37553 12183 37611 12189
rect 38102 12180 38108 12232
rect 38160 12220 38166 12232
rect 38304 12220 38332 12328
rect 39850 12316 39856 12328
rect 39908 12316 39914 12368
rect 39758 12288 39764 12300
rect 38488 12260 39764 12288
rect 38488 12232 38516 12260
rect 39758 12248 39764 12260
rect 39816 12248 39822 12300
rect 40494 12248 40500 12300
rect 40552 12288 40558 12300
rect 40957 12291 41015 12297
rect 40957 12288 40969 12291
rect 40552 12260 40969 12288
rect 40552 12248 40558 12260
rect 40957 12257 40969 12260
rect 41003 12257 41015 12291
rect 40957 12251 41015 12257
rect 38381 12223 38439 12229
rect 38381 12220 38393 12223
rect 38160 12192 38393 12220
rect 38160 12180 38166 12192
rect 38381 12189 38393 12192
rect 38427 12189 38439 12223
rect 38381 12183 38439 12189
rect 38470 12180 38476 12232
rect 38528 12220 38534 12232
rect 38657 12223 38715 12229
rect 38528 12192 38573 12220
rect 38528 12180 38534 12192
rect 38657 12189 38669 12223
rect 38703 12189 38715 12223
rect 38657 12183 38715 12189
rect 34716 12124 35756 12152
rect 38672 12152 38700 12183
rect 38746 12180 38752 12232
rect 38804 12220 38810 12232
rect 39850 12220 39856 12232
rect 38804 12192 38849 12220
rect 39811 12192 39856 12220
rect 38804 12180 38810 12192
rect 39850 12180 39856 12192
rect 39908 12180 39914 12232
rect 40126 12220 40132 12232
rect 40087 12192 40132 12220
rect 40126 12180 40132 12192
rect 40184 12180 40190 12232
rect 41138 12180 41144 12232
rect 41196 12220 41202 12232
rect 41233 12223 41291 12229
rect 41233 12220 41245 12223
rect 41196 12192 41245 12220
rect 41196 12180 41202 12192
rect 41233 12189 41245 12192
rect 41279 12189 41291 12223
rect 41966 12220 41972 12232
rect 41927 12192 41972 12220
rect 41233 12183 41291 12189
rect 41966 12180 41972 12192
rect 42024 12180 42030 12232
rect 43916 12220 43944 12396
rect 46290 12384 46296 12396
rect 46348 12424 46354 12436
rect 46753 12427 46811 12433
rect 46753 12424 46765 12427
rect 46348 12396 46765 12424
rect 46348 12384 46354 12396
rect 46753 12393 46765 12396
rect 46799 12393 46811 12427
rect 46753 12387 46811 12393
rect 47213 12427 47271 12433
rect 47213 12393 47225 12427
rect 47259 12424 47271 12427
rect 48222 12424 48228 12436
rect 47259 12396 48228 12424
rect 47259 12393 47271 12396
rect 47213 12387 47271 12393
rect 48222 12384 48228 12396
rect 48280 12384 48286 12436
rect 49970 12424 49976 12436
rect 48976 12396 49976 12424
rect 43993 12291 44051 12297
rect 43993 12257 44005 12291
rect 44039 12288 44051 12291
rect 47026 12288 47032 12300
rect 44039 12260 47032 12288
rect 44039 12257 44051 12260
rect 43993 12251 44051 12257
rect 47026 12248 47032 12260
rect 47084 12248 47090 12300
rect 48682 12288 48688 12300
rect 48643 12260 48688 12288
rect 48682 12248 48688 12260
rect 48740 12248 48746 12300
rect 48976 12297 49004 12396
rect 49970 12384 49976 12396
rect 50028 12424 50034 12436
rect 50798 12424 50804 12436
rect 50028 12396 50804 12424
rect 50028 12384 50034 12396
rect 50798 12384 50804 12396
rect 50856 12384 50862 12436
rect 51813 12427 51871 12433
rect 51813 12393 51825 12427
rect 51859 12424 51871 12427
rect 51902 12424 51908 12436
rect 51859 12396 51908 12424
rect 51859 12393 51871 12396
rect 51813 12387 51871 12393
rect 51902 12384 51908 12396
rect 51960 12384 51966 12436
rect 53006 12384 53012 12436
rect 53064 12424 53070 12436
rect 53101 12427 53159 12433
rect 53101 12424 53113 12427
rect 53064 12396 53113 12424
rect 53064 12384 53070 12396
rect 53101 12393 53113 12396
rect 53147 12393 53159 12427
rect 53101 12387 53159 12393
rect 53285 12427 53343 12433
rect 53285 12393 53297 12427
rect 53331 12424 53343 12427
rect 54110 12424 54116 12436
rect 53331 12396 54116 12424
rect 53331 12393 53343 12396
rect 53285 12387 53343 12393
rect 54110 12384 54116 12396
rect 54168 12384 54174 12436
rect 54386 12424 54392 12436
rect 54347 12396 54392 12424
rect 54386 12384 54392 12396
rect 54444 12384 54450 12436
rect 49513 12359 49571 12365
rect 49513 12325 49525 12359
rect 49559 12356 49571 12359
rect 49559 12328 51074 12356
rect 49559 12325 49571 12328
rect 49513 12319 49571 12325
rect 48961 12291 49019 12297
rect 48961 12257 48973 12291
rect 49007 12257 49019 12291
rect 49694 12288 49700 12300
rect 48961 12251 49019 12257
rect 49436 12260 49700 12288
rect 49436 12229 49464 12260
rect 49694 12248 49700 12260
rect 49752 12248 49758 12300
rect 51046 12288 51074 12328
rect 51997 12291 52055 12297
rect 51997 12288 52009 12291
rect 51046 12260 52009 12288
rect 51997 12257 52009 12260
rect 52043 12257 52055 12291
rect 51997 12251 52055 12257
rect 53466 12248 53472 12300
rect 53524 12288 53530 12300
rect 54021 12291 54079 12297
rect 54021 12288 54033 12291
rect 53524 12260 54033 12288
rect 53524 12248 53530 12260
rect 54021 12257 54033 12260
rect 54067 12257 54079 12291
rect 54021 12251 54079 12257
rect 54294 12248 54300 12300
rect 54352 12288 54358 12300
rect 54478 12288 54484 12300
rect 54352 12260 54484 12288
rect 54352 12248 54358 12260
rect 54478 12248 54484 12260
rect 54536 12288 54542 12300
rect 57057 12291 57115 12297
rect 57057 12288 57069 12291
rect 54536 12260 57069 12288
rect 54536 12248 54542 12260
rect 57057 12257 57069 12260
rect 57103 12257 57115 12291
rect 57057 12251 57115 12257
rect 44085 12223 44143 12229
rect 44085 12220 44097 12223
rect 43916 12192 44097 12220
rect 44085 12189 44097 12192
rect 44131 12189 44143 12223
rect 44085 12183 44143 12189
rect 45005 12223 45063 12229
rect 45005 12189 45017 12223
rect 45051 12189 45063 12223
rect 45005 12183 45063 12189
rect 49421 12223 49479 12229
rect 49421 12189 49433 12223
rect 49467 12189 49479 12223
rect 49421 12183 49479 12189
rect 49605 12223 49663 12229
rect 49605 12189 49617 12223
rect 49651 12189 49663 12223
rect 50430 12220 50436 12232
rect 50391 12192 50436 12220
rect 49605 12183 49663 12189
rect 39574 12152 39580 12164
rect 38672 12124 39580 12152
rect 39574 12112 39580 12124
rect 39632 12112 39638 12164
rect 39758 12112 39764 12164
rect 39816 12112 39822 12164
rect 42426 12112 42432 12164
rect 42484 12152 42490 12164
rect 42705 12155 42763 12161
rect 42705 12152 42717 12155
rect 42484 12124 42717 12152
rect 42484 12112 42490 12124
rect 42705 12121 42717 12124
rect 42751 12121 42763 12155
rect 42705 12115 42763 12121
rect 43622 12112 43628 12164
rect 43680 12152 43686 12164
rect 45020 12152 45048 12183
rect 43680 12124 45048 12152
rect 45281 12155 45339 12161
rect 43680 12112 43686 12124
rect 45281 12121 45293 12155
rect 45327 12121 45339 12155
rect 45281 12115 45339 12121
rect 17000 12056 17080 12084
rect 17000 12044 17006 12056
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 19426 12084 19432 12096
rect 18288 12056 19432 12084
rect 18288 12044 18294 12056
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 20346 12084 20352 12096
rect 20307 12056 20352 12084
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 23109 12087 23167 12093
rect 23109 12053 23121 12087
rect 23155 12084 23167 12087
rect 23750 12084 23756 12096
rect 23155 12056 23756 12084
rect 23155 12053 23167 12056
rect 23109 12047 23167 12053
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 24394 12044 24400 12096
rect 24452 12084 24458 12096
rect 27614 12084 27620 12096
rect 24452 12056 27620 12084
rect 24452 12044 24458 12056
rect 27614 12044 27620 12056
rect 27672 12044 27678 12096
rect 27709 12087 27767 12093
rect 27709 12053 27721 12087
rect 27755 12084 27767 12087
rect 28258 12084 28264 12096
rect 27755 12056 28264 12084
rect 27755 12053 27767 12056
rect 27709 12047 27767 12053
rect 28258 12044 28264 12056
rect 28316 12044 28322 12096
rect 31481 12087 31539 12093
rect 31481 12053 31493 12087
rect 31527 12084 31539 12087
rect 31570 12084 31576 12096
rect 31527 12056 31576 12084
rect 31527 12053 31539 12056
rect 31481 12047 31539 12053
rect 31570 12044 31576 12056
rect 31628 12044 31634 12096
rect 33134 12044 33140 12096
rect 33192 12084 33198 12096
rect 38286 12084 38292 12096
rect 33192 12056 38292 12084
rect 33192 12044 33198 12056
rect 38286 12044 38292 12056
rect 38344 12044 38350 12096
rect 39776 12084 39804 12112
rect 39945 12087 40003 12093
rect 39945 12084 39957 12087
rect 39776 12056 39957 12084
rect 39945 12053 39957 12056
rect 39991 12053 40003 12087
rect 39945 12047 40003 12053
rect 40034 12044 40040 12096
rect 40092 12084 40098 12096
rect 40313 12087 40371 12093
rect 40313 12084 40325 12087
rect 40092 12056 40325 12084
rect 40092 12044 40098 12056
rect 40313 12053 40325 12056
rect 40359 12053 40371 12087
rect 40313 12047 40371 12053
rect 42150 12044 42156 12096
rect 42208 12084 42214 12096
rect 42797 12087 42855 12093
rect 42797 12084 42809 12087
rect 42208 12056 42809 12084
rect 42208 12044 42214 12056
rect 42797 12053 42809 12056
rect 42843 12084 42855 12087
rect 44174 12084 44180 12096
rect 42843 12056 44180 12084
rect 42843 12053 42855 12056
rect 42797 12047 42855 12053
rect 44174 12044 44180 12056
rect 44232 12044 44238 12096
rect 44453 12087 44511 12093
rect 44453 12053 44465 12087
rect 44499 12084 44511 12087
rect 45296 12084 45324 12115
rect 45370 12112 45376 12164
rect 45428 12152 45434 12164
rect 45428 12124 45770 12152
rect 45428 12112 45434 12124
rect 48222 12112 48228 12164
rect 48280 12112 48286 12164
rect 44499 12056 45324 12084
rect 49620 12084 49648 12183
rect 50430 12180 50436 12192
rect 50488 12180 50494 12232
rect 50709 12223 50767 12229
rect 50709 12189 50721 12223
rect 50755 12189 50767 12223
rect 50709 12183 50767 12189
rect 50724 12152 50752 12183
rect 50798 12180 50804 12232
rect 50856 12220 50862 12232
rect 52089 12223 52147 12229
rect 52089 12220 52101 12223
rect 50856 12192 52101 12220
rect 50856 12180 50862 12192
rect 52089 12189 52101 12192
rect 52135 12189 52147 12223
rect 54205 12223 54263 12229
rect 54205 12220 54217 12223
rect 52089 12183 52147 12189
rect 53484 12192 54217 12220
rect 52546 12152 52552 12164
rect 50724 12124 52552 12152
rect 52546 12112 52552 12124
rect 52604 12152 52610 12164
rect 53374 12152 53380 12164
rect 52604 12124 53380 12152
rect 52604 12112 52610 12124
rect 53374 12112 53380 12124
rect 53432 12112 53438 12164
rect 53484 12161 53512 12192
rect 54205 12189 54217 12192
rect 54251 12220 54263 12223
rect 54251 12192 55214 12220
rect 54251 12189 54263 12192
rect 54205 12183 54263 12189
rect 53469 12155 53527 12161
rect 53469 12121 53481 12155
rect 53515 12121 53527 12155
rect 53469 12115 53527 12121
rect 53834 12112 53840 12164
rect 53892 12152 53898 12164
rect 53929 12155 53987 12161
rect 53929 12152 53941 12155
rect 53892 12124 53941 12152
rect 53892 12112 53898 12124
rect 53929 12121 53941 12124
rect 53975 12121 53987 12155
rect 53929 12115 53987 12121
rect 51074 12084 51080 12096
rect 49620 12056 51080 12084
rect 44499 12053 44511 12056
rect 44453 12047 44511 12053
rect 51074 12044 51080 12056
rect 51132 12044 51138 12096
rect 53006 12044 53012 12096
rect 53064 12084 53070 12096
rect 53259 12087 53317 12093
rect 53259 12084 53271 12087
rect 53064 12056 53271 12084
rect 53064 12044 53070 12056
rect 53259 12053 53271 12056
rect 53305 12053 53317 12087
rect 55186 12084 55214 12192
rect 55674 12180 55680 12232
rect 55732 12180 55738 12232
rect 56778 12152 56784 12164
rect 56739 12124 56784 12152
rect 56778 12112 56784 12124
rect 56836 12112 56842 12164
rect 55306 12084 55312 12096
rect 55186 12056 55312 12084
rect 53259 12047 53317 12053
rect 55306 12044 55312 12056
rect 55364 12044 55370 12096
rect 1104 11994 58880 12016
rect 1104 11942 15398 11994
rect 15450 11942 15462 11994
rect 15514 11942 15526 11994
rect 15578 11942 15590 11994
rect 15642 11942 15654 11994
rect 15706 11942 29846 11994
rect 29898 11942 29910 11994
rect 29962 11942 29974 11994
rect 30026 11942 30038 11994
rect 30090 11942 30102 11994
rect 30154 11942 44294 11994
rect 44346 11942 44358 11994
rect 44410 11942 44422 11994
rect 44474 11942 44486 11994
rect 44538 11942 44550 11994
rect 44602 11942 58880 11994
rect 1104 11920 58880 11942
rect 12250 11880 12256 11892
rect 12211 11852 12256 11880
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 13262 11880 13268 11892
rect 13223 11852 13268 11880
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 14826 11880 14832 11892
rect 14787 11852 14832 11880
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 17586 11840 17592 11892
rect 17644 11880 17650 11892
rect 17865 11883 17923 11889
rect 17865 11880 17877 11883
rect 17644 11852 17877 11880
rect 17644 11840 17650 11852
rect 17865 11849 17877 11852
rect 17911 11849 17923 11883
rect 18690 11880 18696 11892
rect 18651 11852 18696 11880
rect 17865 11843 17923 11849
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 19610 11880 19616 11892
rect 19571 11852 19616 11880
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 23842 11880 23848 11892
rect 22066 11852 23848 11880
rect 11974 11772 11980 11824
rect 12032 11812 12038 11824
rect 13817 11815 13875 11821
rect 13817 11812 13829 11815
rect 12032 11784 13829 11812
rect 12032 11772 12038 11784
rect 13817 11781 13829 11784
rect 13863 11781 13875 11815
rect 13817 11775 13875 11781
rect 16117 11815 16175 11821
rect 16117 11781 16129 11815
rect 16163 11812 16175 11815
rect 16206 11812 16212 11824
rect 16163 11784 16212 11812
rect 16163 11781 16175 11784
rect 16117 11775 16175 11781
rect 16206 11772 16212 11784
rect 16264 11772 16270 11824
rect 16945 11815 17003 11821
rect 16945 11781 16957 11815
rect 16991 11812 17003 11815
rect 19518 11812 19524 11824
rect 16991 11784 19524 11812
rect 16991 11781 17003 11784
rect 16945 11775 17003 11781
rect 19518 11772 19524 11784
rect 19576 11772 19582 11824
rect 22066 11812 22094 11852
rect 23842 11840 23848 11852
rect 23900 11840 23906 11892
rect 24762 11840 24768 11892
rect 24820 11880 24826 11892
rect 25685 11883 25743 11889
rect 25685 11880 25697 11883
rect 24820 11852 25697 11880
rect 24820 11840 24826 11852
rect 25685 11849 25697 11852
rect 25731 11849 25743 11883
rect 25685 11843 25743 11849
rect 26142 11840 26148 11892
rect 26200 11880 26206 11892
rect 26237 11883 26295 11889
rect 26237 11880 26249 11883
rect 26200 11852 26249 11880
rect 26200 11840 26206 11852
rect 26237 11849 26249 11852
rect 26283 11849 26295 11883
rect 30650 11880 30656 11892
rect 30611 11852 30656 11880
rect 26237 11843 26295 11849
rect 30650 11840 30656 11852
rect 30708 11840 30714 11892
rect 30834 11840 30840 11892
rect 30892 11880 30898 11892
rect 31481 11883 31539 11889
rect 31481 11880 31493 11883
rect 30892 11852 31493 11880
rect 30892 11840 30898 11852
rect 31481 11849 31493 11852
rect 31527 11849 31539 11883
rect 33410 11880 33416 11892
rect 33371 11852 33416 11880
rect 31481 11843 31539 11849
rect 33410 11840 33416 11852
rect 33468 11840 33474 11892
rect 33781 11883 33839 11889
rect 33781 11849 33793 11883
rect 33827 11880 33839 11883
rect 34790 11880 34796 11892
rect 33827 11852 34796 11880
rect 33827 11849 33839 11852
rect 33781 11843 33839 11849
rect 34790 11840 34796 11852
rect 34848 11840 34854 11892
rect 35526 11880 35532 11892
rect 35487 11852 35532 11880
rect 35526 11840 35532 11852
rect 35584 11840 35590 11892
rect 35713 11883 35771 11889
rect 35713 11849 35725 11883
rect 35759 11880 35771 11883
rect 38102 11880 38108 11892
rect 35759 11852 38108 11880
rect 35759 11849 35771 11852
rect 35713 11843 35771 11849
rect 38102 11840 38108 11852
rect 38160 11840 38166 11892
rect 40773 11883 40831 11889
rect 40773 11849 40785 11883
rect 40819 11849 40831 11883
rect 40773 11843 40831 11849
rect 23750 11812 23756 11824
rect 19720 11784 22232 11812
rect 23711 11784 23756 11812
rect 12618 11744 12624 11756
rect 12579 11716 12624 11744
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17862 11744 17868 11756
rect 17092 11716 17868 11744
rect 17092 11704 17098 11716
rect 17862 11704 17868 11716
rect 17920 11744 17926 11756
rect 19720 11753 19748 11784
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17920 11716 18613 11744
rect 17920 11704 17926 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 19705 11747 19763 11753
rect 19705 11713 19717 11747
rect 19751 11713 19763 11747
rect 20254 11744 20260 11756
rect 20215 11716 20260 11744
rect 19705 11707 19763 11713
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 21358 11744 21364 11756
rect 20671 11716 21364 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 12713 11679 12771 11685
rect 12713 11645 12725 11679
rect 12759 11676 12771 11679
rect 16850 11676 16856 11688
rect 12759 11648 16856 11676
rect 12759 11645 12771 11648
rect 12713 11639 12771 11645
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 17402 11676 17408 11688
rect 17363 11648 17408 11676
rect 17402 11636 17408 11648
rect 17460 11636 17466 11688
rect 19518 11636 19524 11688
rect 19576 11676 19582 11688
rect 20640 11676 20668 11707
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 21450 11704 21456 11756
rect 21508 11744 21514 11756
rect 22204 11753 22232 11784
rect 23750 11772 23756 11784
rect 23808 11772 23814 11824
rect 27062 11812 27068 11824
rect 24978 11784 27068 11812
rect 27062 11772 27068 11784
rect 27120 11772 27126 11824
rect 28258 11812 28264 11824
rect 28219 11784 28264 11812
rect 28258 11772 28264 11784
rect 28316 11772 28322 11824
rect 29546 11772 29552 11824
rect 29604 11812 29610 11824
rect 30098 11812 30104 11824
rect 29604 11784 30104 11812
rect 29604 11772 29610 11784
rect 30098 11772 30104 11784
rect 30156 11812 30162 11824
rect 30745 11815 30803 11821
rect 30745 11812 30757 11815
rect 30156 11784 30757 11812
rect 30156 11772 30162 11784
rect 30745 11781 30757 11784
rect 30791 11781 30803 11815
rect 35986 11812 35992 11824
rect 30745 11775 30803 11781
rect 31588 11784 35992 11812
rect 31588 11756 31616 11784
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21508 11716 22017 11744
rect 21508 11704 21514 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 23474 11744 23480 11756
rect 23435 11716 23480 11744
rect 22189 11707 22247 11713
rect 23474 11704 23480 11716
rect 23532 11704 23538 11756
rect 30558 11744 30564 11756
rect 30471 11716 30564 11744
rect 30558 11704 30564 11716
rect 30616 11744 30622 11756
rect 31202 11744 31208 11756
rect 30616 11716 31208 11744
rect 30616 11704 30622 11716
rect 31202 11704 31208 11716
rect 31260 11704 31266 11756
rect 31386 11744 31392 11756
rect 31347 11716 31392 11744
rect 31386 11704 31392 11716
rect 31444 11704 31450 11756
rect 31570 11744 31576 11756
rect 31531 11716 31576 11744
rect 31570 11704 31576 11716
rect 31628 11704 31634 11756
rect 31662 11704 31668 11756
rect 31720 11744 31726 11756
rect 32401 11747 32459 11753
rect 32401 11744 32413 11747
rect 31720 11716 32413 11744
rect 31720 11704 31726 11716
rect 32401 11713 32413 11716
rect 32447 11713 32459 11747
rect 32401 11707 32459 11713
rect 32490 11704 32496 11756
rect 32548 11744 32554 11756
rect 32585 11747 32643 11753
rect 32585 11744 32597 11747
rect 32548 11716 32597 11744
rect 32548 11704 32554 11716
rect 32585 11713 32597 11716
rect 32631 11713 32643 11747
rect 33594 11744 33600 11756
rect 33555 11716 33600 11744
rect 32585 11707 32643 11713
rect 33594 11704 33600 11716
rect 33652 11704 33658 11756
rect 33888 11753 33916 11784
rect 35986 11772 35992 11784
rect 36044 11772 36050 11824
rect 37826 11772 37832 11824
rect 37884 11772 37890 11824
rect 38562 11772 38568 11824
rect 38620 11812 38626 11824
rect 40678 11812 40684 11824
rect 38620 11784 39896 11812
rect 38620 11772 38626 11784
rect 33873 11747 33931 11753
rect 33873 11713 33885 11747
rect 33919 11713 33931 11747
rect 34514 11744 34520 11756
rect 34475 11716 34520 11744
rect 33873 11707 33931 11713
rect 34514 11704 34520 11716
rect 34572 11704 34578 11756
rect 34882 11744 34888 11756
rect 34624 11716 34888 11744
rect 19576 11648 20668 11676
rect 21269 11679 21327 11685
rect 19576 11636 19582 11648
rect 21269 11645 21281 11679
rect 21315 11676 21327 11679
rect 22462 11676 22468 11688
rect 21315 11648 22468 11676
rect 21315 11645 21327 11648
rect 21269 11639 21327 11645
rect 22462 11636 22468 11648
rect 22520 11636 22526 11688
rect 23017 11679 23075 11685
rect 23017 11645 23029 11679
rect 23063 11676 23075 11679
rect 24486 11676 24492 11688
rect 23063 11648 24492 11676
rect 23063 11645 23075 11648
rect 23017 11639 23075 11645
rect 24486 11636 24492 11648
rect 24544 11636 24550 11688
rect 27798 11636 27804 11688
rect 27856 11676 27862 11688
rect 28077 11679 28135 11685
rect 28077 11676 28089 11679
rect 27856 11648 28089 11676
rect 27856 11636 27862 11648
rect 28077 11645 28089 11648
rect 28123 11645 28135 11679
rect 28077 11639 28135 11645
rect 28994 11636 29000 11688
rect 29052 11676 29058 11688
rect 29917 11679 29975 11685
rect 29917 11676 29929 11679
rect 29052 11648 29929 11676
rect 29052 11636 29058 11648
rect 29917 11645 29929 11648
rect 29963 11676 29975 11679
rect 30190 11676 30196 11688
rect 29963 11648 30196 11676
rect 29963 11645 29975 11648
rect 29917 11639 29975 11645
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 30377 11679 30435 11685
rect 30377 11645 30389 11679
rect 30423 11676 30435 11679
rect 31110 11676 31116 11688
rect 30423 11648 31116 11676
rect 30423 11645 30435 11648
rect 30377 11639 30435 11645
rect 31110 11636 31116 11648
rect 31168 11676 31174 11688
rect 31168 11648 31754 11676
rect 31168 11636 31174 11648
rect 17678 11608 17684 11620
rect 17639 11580 17684 11608
rect 17678 11568 17684 11580
rect 17736 11568 17742 11620
rect 17788 11580 20944 11608
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 17788 11540 17816 11580
rect 15160 11512 17816 11540
rect 20916 11540 20944 11580
rect 21082 11568 21088 11620
rect 21140 11608 21146 11620
rect 30926 11608 30932 11620
rect 21140 11580 23612 11608
rect 30887 11580 30932 11608
rect 21140 11568 21146 11580
rect 21358 11540 21364 11552
rect 20916 11512 21364 11540
rect 15160 11500 15166 11512
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 23584 11540 23612 11580
rect 30926 11568 30932 11580
rect 30984 11568 30990 11620
rect 31726 11608 31754 11648
rect 32950 11636 32956 11688
rect 33008 11676 33014 11688
rect 34425 11679 34483 11685
rect 34425 11676 34437 11679
rect 33008 11648 34437 11676
rect 33008 11636 33014 11648
rect 34425 11645 34437 11648
rect 34471 11645 34483 11679
rect 34425 11639 34483 11645
rect 34624 11608 34652 11716
rect 34882 11704 34888 11716
rect 34940 11744 34946 11756
rect 35345 11747 35403 11753
rect 35345 11744 35357 11747
rect 34940 11716 35357 11744
rect 34940 11704 34946 11716
rect 35345 11713 35357 11716
rect 35391 11713 35403 11747
rect 35345 11707 35403 11713
rect 35434 11704 35440 11756
rect 35492 11744 35498 11756
rect 35713 11747 35771 11753
rect 35492 11716 35537 11744
rect 35492 11704 35498 11716
rect 35713 11713 35725 11747
rect 35759 11744 35771 11747
rect 35894 11744 35900 11756
rect 35759 11716 35900 11744
rect 35759 11713 35771 11716
rect 35713 11707 35771 11713
rect 35894 11704 35900 11716
rect 35952 11704 35958 11756
rect 36449 11747 36507 11753
rect 36449 11713 36461 11747
rect 36495 11713 36507 11747
rect 36449 11707 36507 11713
rect 31726 11580 34652 11608
rect 25225 11543 25283 11549
rect 25225 11540 25237 11543
rect 23584 11512 25237 11540
rect 25225 11509 25237 11512
rect 25271 11509 25283 11543
rect 25225 11503 25283 11509
rect 32493 11543 32551 11549
rect 32493 11509 32505 11543
rect 32539 11540 32551 11543
rect 32582 11540 32588 11552
rect 32539 11512 32588 11540
rect 32539 11509 32551 11512
rect 32493 11503 32551 11509
rect 32582 11500 32588 11512
rect 32640 11500 32646 11552
rect 34793 11543 34851 11549
rect 34793 11509 34805 11543
rect 34839 11540 34851 11543
rect 35342 11540 35348 11552
rect 34839 11512 35348 11540
rect 34839 11509 34851 11512
rect 34793 11503 34851 11509
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 36262 11540 36268 11552
rect 36223 11512 36268 11540
rect 36262 11500 36268 11512
rect 36320 11500 36326 11552
rect 36464 11540 36492 11707
rect 37369 11679 37427 11685
rect 37369 11645 37381 11679
rect 37415 11676 37427 11679
rect 37642 11676 37648 11688
rect 37415 11648 37648 11676
rect 37415 11645 37427 11648
rect 37369 11639 37427 11645
rect 37642 11636 37648 11648
rect 37700 11676 37706 11688
rect 38470 11676 38476 11688
rect 37700 11648 38476 11676
rect 37700 11636 37706 11648
rect 38470 11636 38476 11648
rect 38528 11636 38534 11688
rect 38838 11676 38844 11688
rect 38799 11648 38844 11676
rect 38838 11636 38844 11648
rect 38896 11636 38902 11688
rect 39117 11679 39175 11685
rect 39117 11645 39129 11679
rect 39163 11645 39175 11679
rect 39574 11676 39580 11688
rect 39535 11648 39580 11676
rect 39117 11639 39175 11645
rect 39132 11608 39160 11639
rect 39574 11636 39580 11648
rect 39632 11636 39638 11688
rect 39868 11685 39896 11784
rect 39960 11784 40684 11812
rect 39960 11753 39988 11784
rect 40678 11772 40684 11784
rect 40736 11772 40742 11824
rect 40788 11812 40816 11843
rect 41966 11840 41972 11892
rect 42024 11880 42030 11892
rect 42613 11883 42671 11889
rect 42613 11880 42625 11883
rect 42024 11852 42625 11880
rect 42024 11840 42030 11852
rect 42613 11849 42625 11852
rect 42659 11849 42671 11883
rect 45370 11880 45376 11892
rect 42613 11843 42671 11849
rect 45112 11852 45376 11880
rect 43625 11815 43683 11821
rect 40788 11784 40908 11812
rect 39945 11747 40003 11753
rect 39945 11713 39957 11747
rect 39991 11713 40003 11747
rect 40586 11744 40592 11756
rect 40547 11716 40592 11744
rect 39945 11707 40003 11713
rect 40586 11704 40592 11716
rect 40644 11704 40650 11756
rect 40773 11747 40831 11753
rect 40773 11713 40785 11747
rect 40819 11713 40831 11747
rect 40773 11707 40831 11713
rect 39853 11679 39911 11685
rect 39853 11645 39865 11679
rect 39899 11645 39911 11679
rect 39853 11639 39911 11645
rect 40218 11608 40224 11620
rect 39132 11580 40224 11608
rect 40218 11568 40224 11580
rect 40276 11568 40282 11620
rect 40788 11608 40816 11707
rect 40880 11676 40908 11784
rect 43625 11781 43637 11815
rect 43671 11812 43683 11815
rect 43806 11812 43812 11824
rect 43671 11784 43812 11812
rect 43671 11781 43683 11784
rect 43625 11775 43683 11781
rect 43806 11772 43812 11784
rect 43864 11772 43870 11824
rect 44174 11772 44180 11824
rect 44232 11812 44238 11824
rect 45112 11812 45140 11852
rect 45370 11840 45376 11852
rect 45428 11840 45434 11892
rect 48314 11880 48320 11892
rect 47964 11852 48320 11880
rect 45186 11812 45192 11824
rect 44232 11784 45192 11812
rect 44232 11772 44238 11784
rect 45186 11772 45192 11784
rect 45244 11772 45250 11824
rect 47964 11821 47992 11852
rect 48314 11840 48320 11852
rect 48372 11880 48378 11892
rect 49510 11880 49516 11892
rect 48372 11852 49516 11880
rect 48372 11840 48378 11852
rect 49510 11840 49516 11852
rect 49568 11840 49574 11892
rect 53926 11880 53932 11892
rect 53887 11852 53932 11880
rect 53926 11840 53932 11852
rect 53984 11840 53990 11892
rect 56597 11883 56655 11889
rect 56597 11849 56609 11883
rect 56643 11880 56655 11883
rect 56778 11880 56784 11892
rect 56643 11852 56784 11880
rect 56643 11849 56655 11852
rect 56597 11843 56655 11849
rect 56778 11840 56784 11852
rect 56836 11840 56842 11892
rect 47949 11815 48007 11821
rect 47949 11781 47961 11815
rect 47995 11781 48007 11815
rect 47949 11775 48007 11781
rect 48222 11772 48228 11824
rect 48280 11812 48286 11824
rect 54205 11815 54263 11821
rect 54205 11812 54217 11815
rect 48280 11784 50200 11812
rect 48280 11772 48286 11784
rect 40954 11704 40960 11756
rect 41012 11744 41018 11756
rect 41417 11747 41475 11753
rect 41417 11744 41429 11747
rect 41012 11716 41429 11744
rect 41012 11704 41018 11716
rect 41417 11713 41429 11716
rect 41463 11713 41475 11747
rect 42426 11744 42432 11756
rect 42387 11716 42432 11744
rect 41417 11707 41475 11713
rect 42426 11704 42432 11716
rect 42484 11704 42490 11756
rect 43714 11704 43720 11756
rect 43772 11744 43778 11756
rect 44453 11747 44511 11753
rect 44453 11744 44465 11747
rect 43772 11716 44465 11744
rect 43772 11704 43778 11716
rect 44453 11713 44465 11716
rect 44499 11713 44511 11747
rect 48130 11744 48136 11756
rect 48091 11716 48136 11744
rect 44453 11707 44511 11713
rect 48130 11704 48136 11716
rect 48188 11704 48194 11756
rect 48777 11747 48835 11753
rect 48777 11744 48789 11747
rect 48332 11716 48789 11744
rect 41325 11679 41383 11685
rect 41325 11676 41337 11679
rect 40880 11648 41337 11676
rect 41325 11645 41337 11648
rect 41371 11645 41383 11679
rect 43438 11676 43444 11688
rect 41325 11639 41383 11645
rect 41524 11648 43444 11676
rect 41524 11608 41552 11648
rect 43438 11636 43444 11648
rect 43496 11636 43502 11688
rect 44729 11679 44787 11685
rect 44729 11645 44741 11679
rect 44775 11676 44787 11679
rect 45094 11676 45100 11688
rect 44775 11648 45100 11676
rect 44775 11645 44787 11648
rect 44729 11639 44787 11645
rect 45094 11636 45100 11648
rect 45152 11636 45158 11688
rect 40788 11580 41552 11608
rect 41616 11580 43760 11608
rect 38194 11540 38200 11552
rect 36464 11512 38200 11540
rect 38194 11500 38200 11512
rect 38252 11500 38258 11552
rect 38286 11500 38292 11552
rect 38344 11540 38350 11552
rect 41616 11540 41644 11580
rect 38344 11512 41644 11540
rect 41693 11543 41751 11549
rect 38344 11500 38350 11512
rect 41693 11509 41705 11543
rect 41739 11540 41751 11543
rect 42426 11540 42432 11552
rect 41739 11512 42432 11540
rect 41739 11509 41751 11512
rect 41693 11503 41751 11509
rect 42426 11500 42432 11512
rect 42484 11500 42490 11552
rect 43732 11549 43760 11580
rect 43717 11543 43775 11549
rect 43717 11509 43729 11543
rect 43763 11540 43775 11543
rect 45370 11540 45376 11552
rect 43763 11512 45376 11540
rect 43763 11509 43775 11512
rect 43717 11503 43775 11509
rect 45370 11500 45376 11512
rect 45428 11500 45434 11552
rect 45462 11500 45468 11552
rect 45520 11540 45526 11552
rect 46201 11543 46259 11549
rect 46201 11540 46213 11543
rect 45520 11512 46213 11540
rect 45520 11500 45526 11512
rect 46201 11509 46213 11512
rect 46247 11509 46259 11543
rect 46201 11503 46259 11509
rect 47854 11500 47860 11552
rect 47912 11540 47918 11552
rect 48332 11549 48360 11716
rect 48777 11713 48789 11716
rect 48823 11713 48835 11747
rect 48777 11707 48835 11713
rect 48961 11747 49019 11753
rect 48961 11713 48973 11747
rect 49007 11744 49019 11747
rect 49694 11744 49700 11756
rect 49007 11716 49700 11744
rect 49007 11713 49019 11716
rect 48961 11707 49019 11713
rect 49694 11704 49700 11716
rect 49752 11704 49758 11756
rect 50172 11753 50200 11784
rect 52932 11784 54217 11812
rect 50157 11747 50215 11753
rect 50157 11713 50169 11747
rect 50203 11744 50215 11747
rect 50890 11744 50896 11756
rect 50203 11716 50896 11744
rect 50203 11713 50215 11716
rect 50157 11707 50215 11713
rect 50890 11704 50896 11716
rect 50948 11704 50954 11756
rect 48498 11636 48504 11688
rect 48556 11676 48562 11688
rect 50430 11676 50436 11688
rect 48556 11648 50436 11676
rect 48556 11636 48562 11648
rect 50430 11636 50436 11648
rect 50488 11676 50494 11688
rect 50801 11679 50859 11685
rect 50801 11676 50813 11679
rect 50488 11648 50813 11676
rect 50488 11636 50494 11648
rect 50801 11645 50813 11648
rect 50847 11645 50859 11679
rect 51074 11676 51080 11688
rect 50987 11648 51080 11676
rect 50801 11639 50859 11645
rect 51074 11636 51080 11648
rect 51132 11676 51138 11688
rect 51994 11676 52000 11688
rect 51132 11648 52000 11676
rect 51132 11636 51138 11648
rect 51994 11636 52000 11648
rect 52052 11636 52058 11688
rect 52932 11685 52960 11784
rect 54205 11781 54217 11784
rect 54251 11812 54263 11815
rect 54251 11784 55168 11812
rect 54251 11781 54263 11784
rect 54205 11775 54263 11781
rect 53101 11747 53159 11753
rect 53101 11713 53113 11747
rect 53147 11744 53159 11747
rect 53282 11744 53288 11756
rect 53147 11716 53288 11744
rect 53147 11713 53159 11716
rect 53101 11707 53159 11713
rect 53282 11704 53288 11716
rect 53340 11704 53346 11756
rect 53926 11744 53932 11756
rect 53887 11716 53932 11744
rect 53926 11704 53932 11716
rect 53984 11704 53990 11756
rect 54021 11747 54079 11753
rect 54021 11713 54033 11747
rect 54067 11744 54079 11747
rect 54110 11744 54116 11756
rect 54067 11716 54116 11744
rect 54067 11713 54079 11716
rect 54021 11707 54079 11713
rect 54110 11704 54116 11716
rect 54168 11744 54174 11756
rect 54938 11744 54944 11756
rect 54168 11716 54944 11744
rect 54168 11704 54174 11716
rect 54938 11704 54944 11716
rect 54996 11704 55002 11756
rect 55140 11744 55168 11784
rect 55306 11744 55312 11756
rect 55140 11716 55312 11744
rect 55306 11704 55312 11716
rect 55364 11744 55370 11756
rect 56229 11747 56287 11753
rect 56229 11744 56241 11747
rect 55364 11716 56241 11744
rect 55364 11704 55370 11716
rect 56229 11713 56241 11716
rect 56275 11713 56287 11747
rect 56229 11707 56287 11713
rect 52917 11679 52975 11685
rect 52917 11645 52929 11679
rect 52963 11645 52975 11679
rect 52917 11639 52975 11645
rect 53006 11636 53012 11688
rect 53064 11676 53070 11688
rect 53064 11648 53157 11676
rect 53064 11636 53070 11648
rect 53190 11636 53196 11688
rect 53248 11676 53254 11688
rect 54849 11679 54907 11685
rect 54849 11676 54861 11679
rect 53248 11648 54861 11676
rect 53248 11636 53254 11648
rect 54849 11645 54861 11648
rect 54895 11645 54907 11679
rect 56134 11676 56140 11688
rect 56095 11648 56140 11676
rect 54849 11639 54907 11645
rect 56134 11636 56140 11648
rect 56192 11636 56198 11688
rect 52638 11568 52644 11620
rect 52696 11608 52702 11620
rect 53024 11608 53052 11636
rect 52696 11580 53052 11608
rect 52696 11568 52702 11580
rect 48317 11543 48375 11549
rect 48317 11540 48329 11543
rect 47912 11512 48329 11540
rect 47912 11500 47918 11512
rect 48317 11509 48329 11512
rect 48363 11509 48375 11543
rect 48317 11503 48375 11509
rect 48958 11500 48964 11552
rect 49016 11540 49022 11552
rect 49145 11543 49203 11549
rect 49145 11540 49157 11543
rect 49016 11512 49157 11540
rect 49016 11500 49022 11512
rect 49145 11509 49157 11512
rect 49191 11509 49203 11543
rect 50246 11540 50252 11552
rect 50207 11512 50252 11540
rect 49145 11503 49203 11509
rect 50246 11500 50252 11512
rect 50304 11500 50310 11552
rect 52086 11540 52092 11552
rect 52047 11512 52092 11540
rect 52086 11500 52092 11512
rect 52144 11500 52150 11552
rect 53098 11500 53104 11552
rect 53156 11540 53162 11552
rect 53469 11543 53527 11549
rect 53469 11540 53481 11543
rect 53156 11512 53481 11540
rect 53156 11500 53162 11512
rect 53469 11509 53481 11512
rect 53515 11509 53527 11543
rect 53469 11503 53527 11509
rect 55217 11543 55275 11549
rect 55217 11509 55229 11543
rect 55263 11540 55275 11543
rect 57790 11540 57796 11552
rect 55263 11512 57796 11540
rect 55263 11509 55275 11512
rect 55217 11503 55275 11509
rect 57790 11500 57796 11512
rect 57848 11500 57854 11552
rect 1104 11450 58880 11472
rect 1104 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 8302 11450
rect 8354 11398 8366 11450
rect 8418 11398 8430 11450
rect 8482 11398 22622 11450
rect 22674 11398 22686 11450
rect 22738 11398 22750 11450
rect 22802 11398 22814 11450
rect 22866 11398 22878 11450
rect 22930 11398 37070 11450
rect 37122 11398 37134 11450
rect 37186 11398 37198 11450
rect 37250 11398 37262 11450
rect 37314 11398 37326 11450
rect 37378 11398 51518 11450
rect 51570 11398 51582 11450
rect 51634 11398 51646 11450
rect 51698 11398 51710 11450
rect 51762 11398 51774 11450
rect 51826 11398 58880 11450
rect 1104 11376 58880 11398
rect 12802 11336 12808 11348
rect 12763 11308 12808 11336
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13412 11308 13553 11336
rect 13412 11296 13418 11308
rect 13541 11305 13553 11308
rect 13587 11336 13599 11339
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13587 11308 14105 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 16666 11336 16672 11348
rect 14093 11299 14151 11305
rect 14568 11308 16672 11336
rect 12253 11271 12311 11277
rect 12253 11237 12265 11271
rect 12299 11268 12311 11271
rect 14568 11268 14596 11308
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 18104 11308 18429 11336
rect 18104 11296 18110 11308
rect 18417 11305 18429 11308
rect 18463 11305 18475 11339
rect 24489 11339 24547 11345
rect 24489 11336 24501 11339
rect 18417 11299 18475 11305
rect 21192 11308 24501 11336
rect 12299 11240 14596 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 16022 11160 16028 11212
rect 16080 11200 16086 11212
rect 19337 11203 19395 11209
rect 19337 11200 19349 11203
rect 16080 11172 19349 11200
rect 16080 11160 16086 11172
rect 19337 11169 19349 11172
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 19702 11160 19708 11212
rect 19760 11200 19766 11212
rect 19886 11200 19892 11212
rect 19760 11172 19892 11200
rect 19760 11160 19766 11172
rect 19886 11160 19892 11172
rect 19944 11160 19950 11212
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11200 20223 11203
rect 20714 11200 20720 11212
rect 20211 11172 20720 11200
rect 20211 11169 20223 11172
rect 20165 11163 20223 11169
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 12161 11135 12219 11141
rect 12161 11132 12173 11135
rect 11940 11104 12173 11132
rect 11940 11092 11946 11104
rect 12161 11101 12173 11104
rect 12207 11101 12219 11135
rect 15102 11132 15108 11144
rect 15063 11104 15108 11132
rect 12161 11095 12219 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 18509 11135 18567 11141
rect 18509 11132 18521 11135
rect 17920 11104 18521 11132
rect 17920 11092 17926 11104
rect 18509 11101 18521 11104
rect 18555 11101 18567 11135
rect 18509 11095 18567 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 19518 11132 19524 11144
rect 19475 11104 19524 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 16022 11064 16028 11076
rect 15983 11036 16028 11064
rect 16022 11024 16028 11036
rect 16080 11024 16086 11076
rect 16574 11024 16580 11076
rect 16632 11024 16638 11076
rect 19720 11064 19748 11160
rect 21192 11132 21220 11308
rect 24489 11305 24501 11308
rect 24535 11305 24547 11339
rect 24489 11299 24547 11305
rect 26973 11339 27031 11345
rect 26973 11305 26985 11339
rect 27019 11336 27031 11339
rect 27338 11336 27344 11348
rect 27019 11308 27344 11336
rect 27019 11305 27031 11308
rect 26973 11299 27031 11305
rect 21358 11228 21364 11280
rect 21416 11268 21422 11280
rect 26988 11268 27016 11299
rect 27338 11296 27344 11308
rect 27396 11296 27402 11348
rect 28626 11336 28632 11348
rect 28587 11308 28632 11336
rect 28626 11296 28632 11308
rect 28684 11296 28690 11348
rect 30926 11296 30932 11348
rect 30984 11336 30990 11348
rect 31573 11339 31631 11345
rect 31573 11336 31585 11339
rect 30984 11308 31585 11336
rect 30984 11296 30990 11308
rect 31573 11305 31585 11308
rect 31619 11336 31631 11339
rect 31662 11336 31668 11348
rect 31619 11308 31668 11336
rect 31619 11305 31631 11308
rect 31573 11299 31631 11305
rect 31662 11296 31668 11308
rect 31720 11296 31726 11348
rect 32950 11336 32956 11348
rect 32911 11308 32956 11336
rect 32950 11296 32956 11308
rect 33008 11296 33014 11348
rect 34514 11296 34520 11348
rect 34572 11336 34578 11348
rect 36817 11339 36875 11345
rect 36817 11336 36829 11339
rect 34572 11308 36829 11336
rect 34572 11296 34578 11308
rect 36817 11305 36829 11308
rect 36863 11305 36875 11339
rect 36817 11299 36875 11305
rect 38657 11339 38715 11345
rect 38657 11305 38669 11339
rect 38703 11336 38715 11339
rect 38838 11336 38844 11348
rect 38703 11308 38844 11336
rect 38703 11305 38715 11308
rect 38657 11299 38715 11305
rect 38838 11296 38844 11308
rect 38896 11296 38902 11348
rect 40405 11339 40463 11345
rect 40405 11305 40417 11339
rect 40451 11336 40463 11339
rect 42702 11336 42708 11348
rect 40451 11308 42708 11336
rect 40451 11305 40463 11308
rect 40405 11299 40463 11305
rect 42702 11296 42708 11308
rect 42760 11296 42766 11348
rect 45094 11336 45100 11348
rect 45055 11308 45100 11336
rect 45094 11296 45100 11308
rect 45152 11296 45158 11348
rect 45370 11296 45376 11348
rect 45428 11336 45434 11348
rect 52086 11336 52092 11348
rect 45428 11308 52092 11336
rect 45428 11296 45434 11308
rect 52086 11296 52092 11308
rect 52144 11336 52150 11348
rect 53190 11336 53196 11348
rect 52144 11308 52408 11336
rect 53151 11308 53196 11336
rect 52144 11296 52150 11308
rect 30558 11268 30564 11280
rect 21416 11240 22140 11268
rect 21416 11228 21422 11240
rect 22112 11209 22140 11240
rect 24596 11240 27016 11268
rect 29748 11240 30564 11268
rect 22097 11203 22155 11209
rect 22097 11169 22109 11203
rect 22143 11169 22155 11203
rect 23842 11200 23848 11212
rect 23803 11172 23848 11200
rect 22097 11163 22155 11169
rect 23842 11160 23848 11172
rect 23900 11160 23906 11212
rect 24394 11132 24400 11144
rect 21192 11104 21298 11132
rect 23506 11104 24400 11132
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 24596 11141 24624 11240
rect 24670 11160 24676 11212
rect 24728 11200 24734 11212
rect 29549 11203 29607 11209
rect 29549 11200 29561 11203
rect 24728 11172 25636 11200
rect 24728 11160 24734 11172
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 24946 11092 24952 11144
rect 25004 11132 25010 11144
rect 25608 11141 25636 11172
rect 28736 11172 29561 11200
rect 28736 11141 28764 11172
rect 29549 11169 29561 11172
rect 29595 11169 29607 11203
rect 29549 11163 29607 11169
rect 29748 11141 29776 11240
rect 30558 11228 30564 11240
rect 30616 11228 30622 11280
rect 40126 11268 40132 11280
rect 36464 11240 40132 11268
rect 30009 11203 30067 11209
rect 30009 11169 30021 11203
rect 30055 11200 30067 11203
rect 30282 11200 30288 11212
rect 30055 11172 30288 11200
rect 30055 11169 30067 11172
rect 30009 11163 30067 11169
rect 30282 11160 30288 11172
rect 30340 11200 30346 11212
rect 30837 11203 30895 11209
rect 30837 11200 30849 11203
rect 30340 11172 30849 11200
rect 30340 11160 30346 11172
rect 30837 11169 30849 11172
rect 30883 11169 30895 11203
rect 35342 11200 35348 11212
rect 35303 11172 35348 11200
rect 30837 11163 30895 11169
rect 35342 11160 35348 11172
rect 35400 11160 35406 11212
rect 35434 11160 35440 11212
rect 35492 11200 35498 11212
rect 36464 11200 36492 11240
rect 40126 11228 40132 11240
rect 40184 11268 40190 11280
rect 40770 11268 40776 11280
rect 40184 11240 40776 11268
rect 40184 11228 40190 11240
rect 40770 11228 40776 11240
rect 40828 11228 40834 11280
rect 40954 11268 40960 11280
rect 40915 11240 40960 11268
rect 40954 11228 40960 11240
rect 41012 11228 41018 11280
rect 43806 11228 43812 11280
rect 43864 11268 43870 11280
rect 48498 11268 48504 11280
rect 43864 11240 48504 11268
rect 43864 11228 43870 11240
rect 48498 11228 48504 11240
rect 48556 11228 48562 11280
rect 49421 11271 49479 11277
rect 49421 11237 49433 11271
rect 49467 11237 49479 11271
rect 49421 11231 49479 11237
rect 35492 11172 36492 11200
rect 35492 11160 35498 11172
rect 36906 11160 36912 11212
rect 36964 11200 36970 11212
rect 37277 11203 37335 11209
rect 37277 11200 37289 11203
rect 36964 11172 37289 11200
rect 36964 11160 36970 11172
rect 37277 11169 37289 11172
rect 37323 11169 37335 11203
rect 37277 11163 37335 11169
rect 39025 11203 39083 11209
rect 39025 11169 39037 11203
rect 39071 11200 39083 11203
rect 39942 11200 39948 11212
rect 39071 11172 39948 11200
rect 39071 11169 39083 11172
rect 39025 11163 39083 11169
rect 39942 11160 39948 11172
rect 40000 11160 40006 11212
rect 40221 11203 40279 11209
rect 40221 11169 40233 11203
rect 40267 11200 40279 11203
rect 40267 11172 41184 11200
rect 40267 11169 40279 11172
rect 40221 11163 40279 11169
rect 25409 11135 25467 11141
rect 25409 11132 25421 11135
rect 25004 11104 25421 11132
rect 25004 11092 25010 11104
rect 25409 11101 25421 11104
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 25593 11135 25651 11141
rect 25593 11101 25605 11135
rect 25639 11101 25651 11135
rect 28537 11135 28595 11141
rect 28537 11132 28549 11135
rect 25593 11095 25651 11101
rect 28184 11104 28549 11132
rect 28184 11076 28212 11104
rect 28537 11101 28549 11104
rect 28583 11101 28595 11135
rect 28537 11095 28595 11101
rect 28721 11135 28779 11141
rect 28721 11101 28733 11135
rect 28767 11101 28779 11135
rect 28721 11095 28779 11101
rect 29733 11135 29791 11141
rect 29733 11101 29745 11135
rect 29779 11101 29791 11135
rect 29733 11095 29791 11101
rect 29825 11135 29883 11141
rect 29825 11101 29837 11135
rect 29871 11101 29883 11135
rect 29825 11095 29883 11101
rect 29917 11135 29975 11141
rect 29917 11101 29929 11135
rect 29963 11132 29975 11135
rect 30374 11132 30380 11144
rect 29963 11104 30380 11132
rect 29963 11101 29975 11104
rect 29917 11095 29975 11101
rect 22370 11064 22376 11076
rect 17880 11036 19748 11064
rect 22331 11036 22376 11064
rect 17880 11008 17908 11036
rect 22370 11024 22376 11036
rect 22428 11024 22434 11076
rect 23842 11024 23848 11076
rect 23900 11064 23906 11076
rect 25498 11064 25504 11076
rect 23900 11036 25504 11064
rect 23900 11024 23906 11036
rect 25498 11024 25504 11036
rect 25556 11024 25562 11076
rect 28077 11067 28135 11073
rect 28077 11033 28089 11067
rect 28123 11064 28135 11067
rect 28166 11064 28172 11076
rect 28123 11036 28172 11064
rect 28123 11033 28135 11036
rect 28077 11027 28135 11033
rect 28166 11024 28172 11036
rect 28224 11024 28230 11076
rect 29840 11064 29868 11095
rect 30374 11092 30380 11104
rect 30432 11092 30438 11144
rect 30745 11135 30803 11141
rect 30745 11101 30757 11135
rect 30791 11101 30803 11135
rect 30745 11095 30803 11101
rect 30929 11135 30987 11141
rect 30929 11101 30941 11135
rect 30975 11132 30987 11135
rect 31018 11132 31024 11144
rect 30975 11104 31024 11132
rect 30975 11101 30987 11104
rect 30929 11095 30987 11101
rect 30098 11064 30104 11076
rect 29840 11036 30104 11064
rect 30098 11024 30104 11036
rect 30156 11064 30162 11076
rect 30760 11064 30788 11095
rect 31018 11092 31024 11104
rect 31076 11132 31082 11144
rect 32493 11135 32551 11141
rect 32493 11132 32505 11135
rect 31076 11104 32505 11132
rect 31076 11092 31082 11104
rect 32493 11101 32505 11104
rect 32539 11101 32551 11135
rect 32493 11095 32551 11101
rect 32582 11092 32588 11144
rect 32640 11132 32646 11144
rect 32769 11135 32827 11141
rect 32640 11104 32685 11132
rect 32640 11092 32646 11104
rect 32769 11101 32781 11135
rect 32815 11101 32827 11135
rect 35066 11132 35072 11144
rect 35027 11104 35072 11132
rect 32769 11095 32827 11101
rect 30156 11036 30788 11064
rect 31481 11067 31539 11073
rect 30156 11024 30162 11036
rect 31481 11033 31493 11067
rect 31527 11064 31539 11067
rect 32784 11064 32812 11095
rect 35066 11092 35072 11104
rect 35124 11092 35130 11144
rect 38102 11132 38108 11144
rect 38063 11104 38108 11132
rect 38102 11092 38108 11104
rect 38160 11092 38166 11144
rect 38470 11092 38476 11144
rect 38528 11132 38534 11144
rect 38933 11135 38991 11141
rect 38933 11132 38945 11135
rect 38528 11104 38945 11132
rect 38528 11092 38534 11104
rect 38933 11101 38945 11104
rect 38979 11101 38991 11135
rect 38933 11095 38991 11101
rect 40034 11092 40040 11144
rect 40092 11132 40098 11144
rect 40129 11135 40187 11141
rect 40129 11132 40141 11135
rect 40092 11104 40141 11132
rect 40092 11092 40098 11104
rect 40129 11101 40141 11104
rect 40175 11101 40187 11135
rect 40129 11095 40187 11101
rect 33505 11067 33563 11073
rect 33505 11064 33517 11067
rect 31527 11036 31708 11064
rect 32784 11036 33517 11064
rect 31527 11033 31539 11036
rect 31481 11027 31539 11033
rect 31680 11008 31708 11036
rect 33505 11033 33517 11036
rect 33551 11064 33563 11067
rect 33594 11064 33600 11076
rect 33551 11036 33600 11064
rect 33551 11033 33563 11036
rect 33505 11027 33563 11033
rect 33594 11024 33600 11036
rect 33652 11064 33658 11076
rect 34057 11067 34115 11073
rect 34057 11064 34069 11067
rect 33652 11036 34069 11064
rect 33652 11024 33658 11036
rect 34057 11033 34069 11036
rect 34103 11064 34115 11067
rect 35434 11064 35440 11076
rect 34103 11036 35440 11064
rect 34103 11033 34115 11036
rect 34057 11027 34115 11033
rect 35434 11024 35440 11036
rect 35492 11024 35498 11076
rect 36630 11064 36636 11076
rect 36543 11036 36636 11064
rect 36630 11024 36636 11036
rect 36688 11064 36694 11076
rect 36688 11036 37136 11064
rect 36688 11024 36694 11036
rect 15197 10999 15255 11005
rect 15197 10965 15209 10999
rect 15243 10996 15255 10999
rect 16206 10996 16212 11008
rect 15243 10968 16212 10996
rect 15243 10965 15255 10968
rect 15197 10959 15255 10965
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 17402 10996 17408 11008
rect 17092 10968 17408 10996
rect 17092 10956 17098 10968
rect 17402 10956 17408 10968
rect 17460 10996 17466 11008
rect 17497 10999 17555 11005
rect 17497 10996 17509 10999
rect 17460 10968 17509 10996
rect 17460 10956 17466 10968
rect 17497 10965 17509 10968
rect 17543 10965 17555 10999
rect 17497 10959 17555 10965
rect 17862 10956 17868 11008
rect 17920 10956 17926 11008
rect 21637 10999 21695 11005
rect 21637 10965 21649 10999
rect 21683 10996 21695 10999
rect 21910 10996 21916 11008
rect 21683 10968 21916 10996
rect 21683 10965 21695 10968
rect 21637 10959 21695 10965
rect 21910 10956 21916 10968
rect 21968 10956 21974 11008
rect 26421 10999 26479 11005
rect 26421 10965 26433 10999
rect 26467 10996 26479 10999
rect 26510 10996 26516 11008
rect 26467 10968 26516 10996
rect 26467 10965 26479 10968
rect 26421 10959 26479 10965
rect 26510 10956 26516 10968
rect 26568 10956 26574 11008
rect 31662 10956 31668 11008
rect 31720 10996 31726 11008
rect 32490 10996 32496 11008
rect 31720 10968 32496 10996
rect 31720 10956 31726 10968
rect 32490 10956 32496 10968
rect 32548 10956 32554 11008
rect 37108 10996 37136 11036
rect 37274 11024 37280 11076
rect 37332 11064 37338 11076
rect 38194 11064 38200 11076
rect 37332 11036 38200 11064
rect 37332 11024 37338 11036
rect 38194 11024 38200 11036
rect 38252 11024 38258 11076
rect 37918 10996 37924 11008
rect 37108 10968 37924 10996
rect 37918 10956 37924 10968
rect 37976 10956 37982 11008
rect 41156 10996 41184 11172
rect 41230 11160 41236 11212
rect 41288 11200 41294 11212
rect 42705 11203 42763 11209
rect 42705 11200 42717 11203
rect 41288 11172 42717 11200
rect 41288 11160 41294 11172
rect 42705 11169 42717 11172
rect 42751 11169 42763 11203
rect 45278 11200 45284 11212
rect 45239 11172 45284 11200
rect 42705 11163 42763 11169
rect 45278 11160 45284 11172
rect 45336 11160 45342 11212
rect 48222 11200 48228 11212
rect 47228 11172 48228 11200
rect 44910 11092 44916 11144
rect 44968 11132 44974 11144
rect 45373 11135 45431 11141
rect 45373 11132 45385 11135
rect 44968 11104 45385 11132
rect 44968 11092 44974 11104
rect 45373 11101 45385 11104
rect 45419 11132 45431 11135
rect 45462 11132 45468 11144
rect 45419 11104 45468 11132
rect 45419 11101 45431 11104
rect 45373 11095 45431 11101
rect 45462 11092 45468 11104
rect 45520 11092 45526 11144
rect 47228 11141 47256 11172
rect 48222 11160 48228 11172
rect 48280 11160 48286 11212
rect 48317 11203 48375 11209
rect 48317 11169 48329 11203
rect 48363 11200 48375 11203
rect 48961 11203 49019 11209
rect 48961 11200 48973 11203
rect 48363 11172 48973 11200
rect 48363 11169 48375 11172
rect 48317 11163 48375 11169
rect 48961 11169 48973 11172
rect 49007 11169 49019 11203
rect 49436 11200 49464 11231
rect 52380 11209 52408 11308
rect 53190 11296 53196 11308
rect 53248 11296 53254 11348
rect 54938 11296 54944 11348
rect 54996 11336 55002 11348
rect 56413 11339 56471 11345
rect 56413 11336 56425 11339
rect 54996 11308 56425 11336
rect 54996 11296 55002 11308
rect 56413 11305 56425 11308
rect 56459 11305 56471 11339
rect 56413 11299 56471 11305
rect 57146 11296 57152 11348
rect 57204 11336 57210 11348
rect 57204 11308 58204 11336
rect 57204 11296 57210 11308
rect 52457 11271 52515 11277
rect 52457 11237 52469 11271
rect 52503 11237 52515 11271
rect 52457 11231 52515 11237
rect 52549 11271 52607 11277
rect 52549 11237 52561 11271
rect 52595 11268 52607 11271
rect 53282 11268 53288 11280
rect 52595 11240 53288 11268
rect 52595 11237 52607 11240
rect 52549 11231 52607 11237
rect 50433 11203 50491 11209
rect 50433 11200 50445 11203
rect 49436 11172 50445 11200
rect 48961 11163 49019 11169
rect 50433 11169 50445 11172
rect 50479 11169 50491 11203
rect 50433 11163 50491 11169
rect 52365 11203 52423 11209
rect 52365 11169 52377 11203
rect 52411 11169 52423 11203
rect 52472 11200 52500 11231
rect 53282 11228 53288 11240
rect 53340 11268 53346 11280
rect 53837 11271 53895 11277
rect 53837 11268 53849 11271
rect 53340 11240 53849 11268
rect 53340 11228 53346 11240
rect 53837 11237 53849 11240
rect 53883 11237 53895 11271
rect 53837 11231 53895 11237
rect 56134 11200 56140 11212
rect 52472 11172 56140 11200
rect 52365 11163 52423 11169
rect 56134 11160 56140 11172
rect 56192 11160 56198 11212
rect 57790 11160 57796 11212
rect 57848 11200 57854 11212
rect 58176 11209 58204 11308
rect 57885 11203 57943 11209
rect 57885 11200 57897 11203
rect 57848 11172 57897 11200
rect 57848 11160 57854 11172
rect 57885 11169 57897 11172
rect 57931 11169 57943 11203
rect 57885 11163 57943 11169
rect 58161 11203 58219 11209
rect 58161 11169 58173 11203
rect 58207 11169 58219 11203
rect 58161 11163 58219 11169
rect 47213 11135 47271 11141
rect 47213 11101 47225 11135
rect 47259 11101 47271 11135
rect 47394 11132 47400 11144
rect 47355 11104 47400 11132
rect 47213 11095 47271 11101
rect 47394 11092 47400 11104
rect 47452 11092 47458 11144
rect 47854 11132 47860 11144
rect 47815 11104 47860 11132
rect 47854 11092 47860 11104
rect 47912 11092 47918 11144
rect 48038 11092 48044 11144
rect 48096 11132 48102 11144
rect 48133 11135 48191 11141
rect 48133 11132 48145 11135
rect 48096 11104 48145 11132
rect 48096 11092 48102 11104
rect 48133 11101 48145 11104
rect 48179 11101 48191 11135
rect 48133 11095 48191 11101
rect 49053 11135 49111 11141
rect 49053 11101 49065 11135
rect 49099 11132 49111 11135
rect 49694 11132 49700 11144
rect 49099 11104 49700 11132
rect 49099 11101 49111 11104
rect 49053 11095 49111 11101
rect 49694 11092 49700 11104
rect 49752 11092 49758 11144
rect 49786 11092 49792 11144
rect 49844 11132 49850 11144
rect 50157 11135 50215 11141
rect 50157 11132 50169 11135
rect 49844 11104 50169 11132
rect 49844 11092 49850 11104
rect 50157 11101 50169 11104
rect 50203 11101 50215 11135
rect 52638 11132 52644 11144
rect 52599 11104 52644 11132
rect 50157 11095 50215 11101
rect 52638 11092 52644 11104
rect 52696 11092 52702 11144
rect 53098 11132 53104 11144
rect 53059 11104 53104 11132
rect 53098 11092 53104 11104
rect 53156 11092 53162 11144
rect 53285 11135 53343 11141
rect 53285 11101 53297 11135
rect 53331 11101 53343 11135
rect 53926 11132 53932 11144
rect 53887 11104 53932 11132
rect 53285 11095 53343 11101
rect 42150 11064 42156 11076
rect 41998 11036 42156 11064
rect 42150 11024 42156 11036
rect 42208 11024 42214 11076
rect 42426 11064 42432 11076
rect 42387 11036 42432 11064
rect 42426 11024 42432 11036
rect 42484 11024 42490 11076
rect 47305 11067 47363 11073
rect 47305 11033 47317 11067
rect 47351 11064 47363 11067
rect 47949 11067 48007 11073
rect 47949 11064 47961 11067
rect 47351 11036 47961 11064
rect 47351 11033 47363 11036
rect 47305 11027 47363 11033
rect 47949 11033 47961 11036
rect 47995 11033 48007 11067
rect 47949 11027 48007 11033
rect 50890 11024 50896 11076
rect 50948 11024 50954 11076
rect 51994 11024 52000 11076
rect 52052 11064 52058 11076
rect 53300 11064 53328 11095
rect 53926 11092 53932 11104
rect 53984 11092 53990 11144
rect 52052 11036 53328 11064
rect 52052 11024 52058 11036
rect 56594 11024 56600 11076
rect 56652 11064 56658 11076
rect 56652 11036 56718 11064
rect 56652 11024 56658 11036
rect 42334 10996 42340 11008
rect 41156 10968 42340 10996
rect 42334 10956 42340 10968
rect 42392 10956 42398 11008
rect 43530 10996 43536 11008
rect 43491 10968 43536 10996
rect 43530 10956 43536 10968
rect 43588 10956 43594 11008
rect 47394 10956 47400 11008
rect 47452 10996 47458 11008
rect 48130 10996 48136 11008
rect 47452 10968 48136 10996
rect 47452 10956 47458 10968
rect 48130 10956 48136 10968
rect 48188 10956 48194 11008
rect 51902 10996 51908 11008
rect 51863 10968 51908 10996
rect 51902 10956 51908 10968
rect 51960 10956 51966 11008
rect 1104 10906 58880 10928
rect 1104 10854 15398 10906
rect 15450 10854 15462 10906
rect 15514 10854 15526 10906
rect 15578 10854 15590 10906
rect 15642 10854 15654 10906
rect 15706 10854 29846 10906
rect 29898 10854 29910 10906
rect 29962 10854 29974 10906
rect 30026 10854 30038 10906
rect 30090 10854 30102 10906
rect 30154 10854 44294 10906
rect 44346 10854 44358 10906
rect 44410 10854 44422 10906
rect 44474 10854 44486 10906
rect 44538 10854 44550 10906
rect 44602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1912 10764 1961 10792
rect 1912 10752 1918 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 1949 10755 2007 10761
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16117 10795 16175 10801
rect 16117 10792 16129 10795
rect 16080 10764 16129 10792
rect 16080 10752 16086 10764
rect 16117 10761 16129 10764
rect 16163 10761 16175 10795
rect 16117 10755 16175 10761
rect 17129 10795 17187 10801
rect 17129 10761 17141 10795
rect 17175 10792 17187 10795
rect 17954 10792 17960 10804
rect 17175 10764 17960 10792
rect 17175 10761 17187 10764
rect 17129 10755 17187 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 18598 10752 18604 10804
rect 18656 10792 18662 10804
rect 21174 10792 21180 10804
rect 18656 10764 20760 10792
rect 21135 10764 21180 10792
rect 18656 10752 18662 10764
rect 16574 10724 16580 10736
rect 15870 10696 16580 10724
rect 16574 10684 16580 10696
rect 16632 10724 16638 10736
rect 17586 10724 17592 10736
rect 16632 10696 17592 10724
rect 16632 10684 16638 10696
rect 17586 10684 17592 10696
rect 17644 10684 17650 10736
rect 17681 10727 17739 10733
rect 17681 10693 17693 10727
rect 17727 10724 17739 10727
rect 17862 10724 17868 10736
rect 17727 10696 17868 10724
rect 17727 10693 17739 10696
rect 17681 10687 17739 10693
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1857 10659 1915 10665
rect 1857 10656 1869 10659
rect 1636 10628 1869 10656
rect 1636 10616 1642 10628
rect 1857 10625 1869 10628
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 17696 10656 17724 10687
rect 17862 10684 17868 10696
rect 17920 10684 17926 10736
rect 20438 10724 20444 10736
rect 20399 10696 20444 10724
rect 20438 10684 20444 10696
rect 20496 10684 20502 10736
rect 16264 10628 17724 10656
rect 16264 10616 16270 10628
rect 19334 10616 19340 10668
rect 19392 10616 19398 10668
rect 20732 10665 20760 10764
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 21910 10752 21916 10804
rect 21968 10792 21974 10804
rect 26421 10795 26479 10801
rect 21968 10764 25452 10792
rect 21968 10752 21974 10764
rect 22189 10727 22247 10733
rect 22189 10693 22201 10727
rect 22235 10724 22247 10727
rect 22370 10724 22376 10736
rect 22235 10696 22376 10724
rect 22235 10693 22247 10696
rect 22189 10687 22247 10693
rect 22370 10684 22376 10696
rect 22428 10684 22434 10736
rect 24486 10684 24492 10736
rect 24544 10724 24550 10736
rect 24581 10727 24639 10733
rect 24581 10724 24593 10727
rect 24544 10696 24593 10724
rect 24544 10684 24550 10696
rect 24581 10693 24593 10696
rect 24627 10693 24639 10727
rect 24581 10687 24639 10693
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10656 20775 10659
rect 21174 10656 21180 10668
rect 20763 10628 21180 10656
rect 20763 10625 20775 10628
rect 20717 10619 20775 10625
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 21910 10656 21916 10668
rect 21871 10628 21916 10656
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 25424 10665 25452 10764
rect 26421 10761 26433 10795
rect 26467 10792 26479 10795
rect 36357 10795 36415 10801
rect 26467 10764 32628 10792
rect 26467 10761 26479 10764
rect 26421 10755 26479 10761
rect 29086 10724 29092 10736
rect 26988 10696 29092 10724
rect 25409 10659 25467 10665
rect 25409 10625 25421 10659
rect 25455 10625 25467 10659
rect 25409 10619 25467 10625
rect 25498 10616 25504 10668
rect 25556 10656 25562 10668
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 25556 10628 25605 10656
rect 25556 10616 25562 10628
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 25593 10619 25651 10625
rect 14369 10591 14427 10597
rect 14369 10588 14381 10591
rect 13832 10560 14381 10588
rect 13832 10464 13860 10560
rect 14369 10557 14381 10560
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 16669 10591 16727 10597
rect 16669 10588 16681 10591
rect 14691 10560 16681 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 16669 10557 16681 10560
rect 16715 10588 16727 10591
rect 17678 10588 17684 10600
rect 16715 10560 17684 10588
rect 16715 10557 16727 10560
rect 16669 10551 16727 10557
rect 17678 10548 17684 10560
rect 17736 10588 17742 10600
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 17736 10560 18981 10588
rect 17736 10548 17742 10560
rect 18969 10557 18981 10560
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 20346 10548 20352 10600
rect 20404 10588 20410 10600
rect 20404 10560 20668 10588
rect 20404 10548 20410 10560
rect 17034 10520 17040 10532
rect 16995 10492 17040 10520
rect 17034 10480 17040 10492
rect 17092 10480 17098 10532
rect 20640 10520 20668 10560
rect 23566 10548 23572 10600
rect 23624 10588 23630 10600
rect 24305 10591 24363 10597
rect 24305 10588 24317 10591
rect 23624 10560 24317 10588
rect 23624 10548 23630 10560
rect 24305 10557 24317 10560
rect 24351 10588 24363 10591
rect 24486 10588 24492 10600
rect 24351 10560 24492 10588
rect 24351 10557 24363 10560
rect 24305 10551 24363 10557
rect 24486 10548 24492 10560
rect 24544 10548 24550 10600
rect 24765 10591 24823 10597
rect 24765 10557 24777 10591
rect 24811 10588 24823 10591
rect 26988 10588 27016 10696
rect 29086 10684 29092 10696
rect 29144 10684 29150 10736
rect 29178 10684 29184 10736
rect 29236 10724 29242 10736
rect 29733 10727 29791 10733
rect 29733 10724 29745 10727
rect 29236 10696 29745 10724
rect 29236 10684 29242 10696
rect 29733 10693 29745 10696
rect 29779 10693 29791 10727
rect 29733 10687 29791 10693
rect 31754 10616 31760 10668
rect 31812 10656 31818 10668
rect 32309 10659 32367 10665
rect 32309 10656 32321 10659
rect 31812 10628 32321 10656
rect 31812 10616 31818 10628
rect 32309 10625 32321 10628
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 27154 10588 27160 10600
rect 24811 10560 27016 10588
rect 27115 10560 27160 10588
rect 24811 10557 24823 10560
rect 24765 10551 24823 10557
rect 27154 10548 27160 10560
rect 27212 10548 27218 10600
rect 28629 10591 28687 10597
rect 28629 10557 28641 10591
rect 28675 10557 28687 10591
rect 28629 10551 28687 10557
rect 28813 10591 28871 10597
rect 28813 10557 28825 10591
rect 28859 10557 28871 10591
rect 29546 10588 29552 10600
rect 29507 10560 29552 10588
rect 28813 10551 28871 10557
rect 28644 10520 28672 10551
rect 20640 10492 28672 10520
rect 28828 10520 28856 10551
rect 29546 10548 29552 10560
rect 29604 10548 29610 10600
rect 30190 10548 30196 10600
rect 30248 10588 30254 10600
rect 30742 10588 30748 10600
rect 30248 10560 30748 10588
rect 30248 10548 30254 10560
rect 30742 10548 30748 10560
rect 30800 10548 30806 10600
rect 32217 10591 32275 10597
rect 32217 10588 32229 10591
rect 31726 10560 32229 10588
rect 30374 10520 30380 10532
rect 28828 10492 30380 10520
rect 30374 10480 30380 10492
rect 30432 10480 30438 10532
rect 30650 10480 30656 10532
rect 30708 10520 30714 10532
rect 31726 10520 31754 10560
rect 32217 10557 32229 10560
rect 32263 10557 32275 10591
rect 32217 10551 32275 10557
rect 30708 10492 31754 10520
rect 32600 10520 32628 10764
rect 36357 10761 36369 10795
rect 36403 10792 36415 10795
rect 36630 10792 36636 10804
rect 36403 10764 36636 10792
rect 36403 10761 36415 10764
rect 36357 10755 36415 10761
rect 36630 10752 36636 10764
rect 36688 10752 36694 10804
rect 38470 10752 38476 10804
rect 38528 10792 38534 10804
rect 40954 10792 40960 10804
rect 38528 10764 40960 10792
rect 38528 10752 38534 10764
rect 40954 10752 40960 10764
rect 41012 10752 41018 10804
rect 42334 10752 42340 10804
rect 42392 10792 42398 10804
rect 42429 10795 42487 10801
rect 42429 10792 42441 10795
rect 42392 10764 42441 10792
rect 42392 10752 42398 10764
rect 42429 10761 42441 10764
rect 42475 10761 42487 10795
rect 42429 10755 42487 10761
rect 43257 10795 43315 10801
rect 43257 10761 43269 10795
rect 43303 10792 43315 10795
rect 43438 10792 43444 10804
rect 43303 10764 43444 10792
rect 43303 10761 43315 10764
rect 43257 10755 43315 10761
rect 43438 10752 43444 10764
rect 43496 10752 43502 10804
rect 48869 10795 48927 10801
rect 48869 10761 48881 10795
rect 48915 10792 48927 10795
rect 49421 10795 49479 10801
rect 49421 10792 49433 10795
rect 48915 10764 49433 10792
rect 48915 10761 48927 10764
rect 48869 10755 48927 10761
rect 49421 10761 49433 10764
rect 49467 10761 49479 10795
rect 49421 10755 49479 10761
rect 51997 10795 52055 10801
rect 51997 10761 52009 10795
rect 52043 10792 52055 10795
rect 52638 10792 52644 10804
rect 52043 10764 52644 10792
rect 52043 10761 52055 10764
rect 51997 10755 52055 10761
rect 52638 10752 52644 10764
rect 52696 10752 52702 10804
rect 33778 10724 33784 10736
rect 33739 10696 33784 10724
rect 33778 10684 33784 10696
rect 33836 10684 33842 10736
rect 35529 10727 35587 10733
rect 35529 10693 35541 10727
rect 35575 10724 35587 10727
rect 38930 10724 38936 10736
rect 35575 10696 38936 10724
rect 35575 10693 35587 10696
rect 35529 10687 35587 10693
rect 38930 10684 38936 10696
rect 38988 10724 38994 10736
rect 39025 10727 39083 10733
rect 39025 10724 39037 10727
rect 38988 10696 39037 10724
rect 38988 10684 38994 10696
rect 39025 10693 39037 10696
rect 39071 10693 39083 10727
rect 39025 10687 39083 10693
rect 39206 10684 39212 10736
rect 39264 10724 39270 10736
rect 41233 10727 41291 10733
rect 41233 10724 41245 10727
rect 39264 10696 41245 10724
rect 39264 10684 39270 10696
rect 41233 10693 41245 10696
rect 41279 10693 41291 10727
rect 41233 10687 41291 10693
rect 41417 10727 41475 10733
rect 41417 10693 41429 10727
rect 41463 10724 41475 10727
rect 41463 10696 42840 10724
rect 41463 10693 41475 10696
rect 41417 10687 41475 10693
rect 36541 10659 36599 10665
rect 36541 10625 36553 10659
rect 36587 10656 36599 10659
rect 37274 10656 37280 10668
rect 36587 10628 37280 10656
rect 36587 10625 36599 10628
rect 36541 10619 36599 10625
rect 37274 10616 37280 10628
rect 37332 10616 37338 10668
rect 37734 10656 37740 10668
rect 37695 10628 37740 10656
rect 37734 10616 37740 10628
rect 37792 10616 37798 10668
rect 37829 10659 37887 10665
rect 37829 10625 37841 10659
rect 37875 10625 37887 10659
rect 37829 10619 37887 10625
rect 37553 10591 37611 10597
rect 37553 10557 37565 10591
rect 37599 10557 37611 10591
rect 37844 10588 37872 10619
rect 37918 10616 37924 10668
rect 37976 10656 37982 10668
rect 38381 10659 38439 10665
rect 38381 10656 38393 10659
rect 37976 10628 38393 10656
rect 37976 10616 37982 10628
rect 38381 10625 38393 10628
rect 38427 10625 38439 10659
rect 40310 10656 40316 10668
rect 38381 10619 38439 10625
rect 38488 10628 40316 10656
rect 38488 10588 38516 10628
rect 40310 10616 40316 10628
rect 40368 10616 40374 10668
rect 42518 10656 42524 10668
rect 41984 10628 42524 10656
rect 37844 10560 38516 10588
rect 38565 10591 38623 10597
rect 37553 10551 37611 10557
rect 38565 10557 38577 10591
rect 38611 10588 38623 10591
rect 41984 10588 42012 10628
rect 42518 10616 42524 10628
rect 42576 10616 42582 10668
rect 42610 10616 42616 10668
rect 42668 10656 42674 10668
rect 42705 10659 42763 10665
rect 42705 10656 42717 10659
rect 42668 10628 42717 10656
rect 42668 10616 42674 10628
rect 42705 10625 42717 10628
rect 42751 10625 42763 10659
rect 42705 10619 42763 10625
rect 38611 10560 42012 10588
rect 42429 10591 42487 10597
rect 38611 10557 38623 10560
rect 38565 10551 38623 10557
rect 42429 10557 42441 10591
rect 42475 10588 42487 10591
rect 42812 10588 42840 10696
rect 48038 10684 48044 10736
rect 48096 10724 48102 10736
rect 49694 10724 49700 10736
rect 48096 10696 48728 10724
rect 49607 10696 49700 10724
rect 48096 10684 48102 10696
rect 43349 10659 43407 10665
rect 43349 10625 43361 10659
rect 43395 10656 43407 10659
rect 43530 10656 43536 10668
rect 43395 10628 43536 10656
rect 43395 10625 43407 10628
rect 43349 10619 43407 10625
rect 43530 10616 43536 10628
rect 43588 10616 43594 10668
rect 43806 10616 43812 10668
rect 43864 10656 43870 10668
rect 48700 10665 48728 10696
rect 49694 10684 49700 10696
rect 49752 10724 49758 10736
rect 51721 10727 51779 10733
rect 51721 10724 51733 10727
rect 49752 10696 51733 10724
rect 49752 10684 49758 10696
rect 51721 10693 51733 10696
rect 51767 10724 51779 10727
rect 51902 10724 51908 10736
rect 51767 10696 51908 10724
rect 51767 10693 51779 10696
rect 51721 10687 51779 10693
rect 51902 10684 51908 10696
rect 51960 10684 51966 10736
rect 44269 10659 44327 10665
rect 44269 10656 44281 10659
rect 43864 10628 44281 10656
rect 43864 10616 43870 10628
rect 44269 10625 44281 10628
rect 44315 10625 44327 10659
rect 44269 10619 44327 10625
rect 48685 10659 48743 10665
rect 48685 10625 48697 10659
rect 48731 10625 48743 10659
rect 48958 10656 48964 10668
rect 48919 10628 48964 10656
rect 48685 10619 48743 10625
rect 48958 10616 48964 10628
rect 49016 10616 49022 10668
rect 49421 10659 49479 10665
rect 49421 10625 49433 10659
rect 49467 10625 49479 10659
rect 49421 10619 49479 10625
rect 43824 10588 43852 10616
rect 42475 10560 43852 10588
rect 43993 10591 44051 10597
rect 42475 10557 42487 10560
rect 42429 10551 42487 10557
rect 43993 10557 44005 10591
rect 44039 10557 44051 10591
rect 43993 10551 44051 10557
rect 37458 10520 37464 10532
rect 32600 10492 37464 10520
rect 30708 10480 30714 10492
rect 37458 10480 37464 10492
rect 37516 10480 37522 10532
rect 37568 10520 37596 10551
rect 40034 10520 40040 10532
rect 37568 10492 40040 10520
rect 40034 10480 40040 10492
rect 40092 10480 40098 10532
rect 41138 10480 41144 10532
rect 41196 10520 41202 10532
rect 42613 10523 42671 10529
rect 42613 10520 42625 10523
rect 41196 10492 42625 10520
rect 41196 10480 41202 10492
rect 42613 10489 42625 10492
rect 42659 10489 42671 10523
rect 42613 10483 42671 10489
rect 13814 10452 13820 10464
rect 13775 10424 13820 10452
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 20990 10452 20996 10464
rect 18555 10424 20996 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 32582 10452 32588 10464
rect 32543 10424 32588 10452
rect 32582 10412 32588 10424
rect 32640 10412 32646 10464
rect 37829 10455 37887 10461
rect 37829 10421 37841 10455
rect 37875 10452 37887 10455
rect 39942 10452 39948 10464
rect 37875 10424 39948 10452
rect 37875 10421 37887 10424
rect 37829 10415 37887 10421
rect 39942 10412 39948 10424
rect 40000 10412 40006 10464
rect 40218 10412 40224 10464
rect 40276 10452 40282 10464
rect 40313 10455 40371 10461
rect 40313 10452 40325 10455
rect 40276 10424 40325 10452
rect 40276 10412 40282 10424
rect 40313 10421 40325 10424
rect 40359 10421 40371 10455
rect 40313 10415 40371 10421
rect 43530 10412 43536 10464
rect 43588 10452 43594 10464
rect 44008 10452 44036 10551
rect 48130 10548 48136 10600
rect 48188 10588 48194 10600
rect 49436 10588 49464 10619
rect 49510 10616 49516 10668
rect 49568 10656 49574 10668
rect 51350 10656 51356 10668
rect 49568 10628 51356 10656
rect 49568 10616 49574 10628
rect 51350 10616 51356 10628
rect 51408 10656 51414 10668
rect 51629 10659 51687 10665
rect 51629 10656 51641 10659
rect 51408 10628 51641 10656
rect 51408 10616 51414 10628
rect 51629 10625 51641 10628
rect 51675 10625 51687 10659
rect 51629 10619 51687 10625
rect 51813 10659 51871 10665
rect 51813 10625 51825 10659
rect 51859 10656 51871 10659
rect 52362 10656 52368 10668
rect 51859 10628 52368 10656
rect 51859 10625 51871 10628
rect 51813 10619 51871 10625
rect 52362 10616 52368 10628
rect 52420 10656 52426 10668
rect 53009 10659 53067 10665
rect 53009 10656 53021 10659
rect 52420 10628 53021 10656
rect 52420 10616 52426 10628
rect 53009 10625 53021 10628
rect 53055 10656 53067 10659
rect 56042 10656 56048 10668
rect 53055 10628 56048 10656
rect 53055 10625 53067 10628
rect 53009 10619 53067 10625
rect 56042 10616 56048 10628
rect 56100 10616 56106 10668
rect 52917 10591 52975 10597
rect 52917 10588 52929 10591
rect 48188 10560 51074 10588
rect 48188 10548 48194 10560
rect 48501 10523 48559 10529
rect 48501 10489 48513 10523
rect 48547 10520 48559 10523
rect 51046 10520 51074 10560
rect 51552 10560 52929 10588
rect 51442 10520 51448 10532
rect 48547 10492 49832 10520
rect 51046 10492 51448 10520
rect 48547 10489 48559 10492
rect 48501 10483 48559 10489
rect 45370 10452 45376 10464
rect 43588 10424 45376 10452
rect 43588 10412 43594 10424
rect 45370 10412 45376 10424
rect 45428 10412 45434 10464
rect 45554 10412 45560 10464
rect 45612 10452 45618 10464
rect 47673 10455 47731 10461
rect 47673 10452 47685 10455
rect 45612 10424 47685 10452
rect 45612 10412 45618 10424
rect 47673 10421 47685 10424
rect 47719 10452 47731 10455
rect 48038 10452 48044 10464
rect 47719 10424 48044 10452
rect 47719 10421 47731 10424
rect 47673 10415 47731 10421
rect 48038 10412 48044 10424
rect 48096 10412 48102 10464
rect 49804 10452 49832 10492
rect 51442 10480 51448 10492
rect 51500 10480 51506 10532
rect 51552 10452 51580 10560
rect 52917 10557 52929 10560
rect 52963 10557 52975 10591
rect 52917 10551 52975 10557
rect 53377 10523 53435 10529
rect 53377 10489 53389 10523
rect 53423 10520 53435 10523
rect 54570 10520 54576 10532
rect 53423 10492 54576 10520
rect 53423 10489 53435 10492
rect 53377 10483 53435 10489
rect 54570 10480 54576 10492
rect 54628 10480 54634 10532
rect 49804 10424 51580 10452
rect 1104 10362 58880 10384
rect 1104 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 8302 10362
rect 8354 10310 8366 10362
rect 8418 10310 8430 10362
rect 8482 10310 22622 10362
rect 22674 10310 22686 10362
rect 22738 10310 22750 10362
rect 22802 10310 22814 10362
rect 22866 10310 22878 10362
rect 22930 10310 37070 10362
rect 37122 10310 37134 10362
rect 37186 10310 37198 10362
rect 37250 10310 37262 10362
rect 37314 10310 37326 10362
rect 37378 10310 51518 10362
rect 51570 10310 51582 10362
rect 51634 10310 51646 10362
rect 51698 10310 51710 10362
rect 51762 10310 51774 10362
rect 51826 10310 58880 10362
rect 1104 10288 58880 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 16206 10248 16212 10260
rect 16167 10220 16212 10248
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 19613 10251 19671 10257
rect 19613 10217 19625 10251
rect 19659 10248 19671 10251
rect 24578 10248 24584 10260
rect 19659 10220 24584 10248
rect 19659 10217 19671 10220
rect 19613 10211 19671 10217
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 30466 10248 30472 10260
rect 25884 10220 30472 10248
rect 16666 10140 16672 10192
rect 16724 10180 16730 10192
rect 21085 10183 21143 10189
rect 21085 10180 21097 10183
rect 16724 10152 21097 10180
rect 16724 10140 16730 10152
rect 21085 10149 21097 10152
rect 21131 10149 21143 10183
rect 21085 10143 21143 10149
rect 21174 10140 21180 10192
rect 21232 10180 21238 10192
rect 25884 10180 25912 10220
rect 30466 10208 30472 10220
rect 30524 10208 30530 10260
rect 30650 10248 30656 10260
rect 30611 10220 30656 10248
rect 30650 10208 30656 10220
rect 30708 10208 30714 10260
rect 31018 10208 31024 10260
rect 31076 10248 31082 10260
rect 31205 10251 31263 10257
rect 31205 10248 31217 10251
rect 31076 10220 31217 10248
rect 31076 10208 31082 10220
rect 31205 10217 31217 10220
rect 31251 10217 31263 10251
rect 31478 10248 31484 10260
rect 31439 10220 31484 10248
rect 31205 10211 31263 10217
rect 31478 10208 31484 10220
rect 31536 10248 31542 10260
rect 31536 10220 32444 10248
rect 31536 10208 31542 10220
rect 27706 10180 27712 10192
rect 21232 10152 25912 10180
rect 26988 10152 27712 10180
rect 21232 10140 21238 10152
rect 18138 10112 18144 10124
rect 18051 10084 18144 10112
rect 18138 10072 18144 10084
rect 18196 10112 18202 10124
rect 23845 10115 23903 10121
rect 18196 10084 20484 10112
rect 18196 10072 18202 10084
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10044 19579 10047
rect 20254 10044 20260 10056
rect 19567 10016 20260 10044
rect 19567 10013 19579 10016
rect 19521 10007 19579 10013
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 20349 9979 20407 9985
rect 20349 9976 20361 9979
rect 19392 9948 20361 9976
rect 19392 9936 19398 9948
rect 20349 9945 20361 9948
rect 20395 9945 20407 9979
rect 20456 9976 20484 10084
rect 23845 10081 23857 10115
rect 23891 10112 23903 10115
rect 26234 10112 26240 10124
rect 23891 10084 26240 10112
rect 23891 10081 23903 10084
rect 23845 10075 23903 10081
rect 26234 10072 26240 10084
rect 26292 10072 26298 10124
rect 26510 10112 26516 10124
rect 26471 10084 26516 10112
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 26697 10115 26755 10121
rect 26697 10081 26709 10115
rect 26743 10112 26755 10115
rect 26988 10112 27016 10152
rect 27706 10140 27712 10152
rect 27764 10140 27770 10192
rect 28258 10140 28264 10192
rect 28316 10180 28322 10192
rect 28316 10152 29040 10180
rect 28316 10140 28322 10152
rect 27154 10112 27160 10124
rect 26743 10084 27016 10112
rect 27115 10084 27160 10112
rect 26743 10081 26755 10084
rect 26697 10075 26755 10081
rect 27154 10072 27160 10084
rect 27212 10072 27218 10124
rect 28718 10072 28724 10124
rect 28776 10112 28782 10124
rect 29012 10121 29040 10152
rect 29362 10140 29368 10192
rect 29420 10180 29426 10192
rect 29825 10183 29883 10189
rect 29825 10180 29837 10183
rect 29420 10152 29837 10180
rect 29420 10140 29426 10152
rect 29825 10149 29837 10152
rect 29871 10149 29883 10183
rect 31662 10180 31668 10192
rect 29825 10143 29883 10149
rect 31496 10152 31668 10180
rect 28813 10115 28871 10121
rect 28813 10112 28825 10115
rect 28776 10084 28825 10112
rect 28776 10072 28782 10084
rect 28813 10081 28825 10084
rect 28859 10081 28871 10115
rect 28813 10075 28871 10081
rect 28997 10115 29055 10121
rect 28997 10081 29009 10115
rect 29043 10081 29055 10115
rect 28997 10075 29055 10081
rect 30009 10115 30067 10121
rect 30009 10081 30021 10115
rect 30055 10112 30067 10115
rect 30561 10115 30619 10121
rect 30561 10112 30573 10115
rect 30055 10084 30573 10112
rect 30055 10081 30067 10084
rect 30009 10075 30067 10081
rect 30561 10081 30573 10084
rect 30607 10081 30619 10115
rect 30561 10075 30619 10081
rect 30745 10115 30803 10121
rect 30745 10081 30757 10115
rect 30791 10112 30803 10115
rect 30834 10112 30840 10124
rect 30791 10084 30840 10112
rect 30791 10081 30803 10084
rect 30745 10075 30803 10081
rect 30834 10072 30840 10084
rect 30892 10072 30898 10124
rect 31496 10121 31524 10152
rect 31662 10140 31668 10152
rect 31720 10140 31726 10192
rect 32416 10180 32444 10220
rect 32582 10208 32588 10260
rect 32640 10248 32646 10260
rect 34958 10251 35016 10257
rect 34958 10248 34970 10251
rect 32640 10220 34970 10248
rect 32640 10208 32646 10220
rect 34958 10217 34970 10220
rect 35004 10217 35016 10251
rect 40586 10248 40592 10260
rect 40547 10220 40592 10248
rect 34958 10211 35016 10217
rect 40586 10208 40592 10220
rect 40644 10208 40650 10260
rect 40770 10208 40776 10260
rect 40828 10248 40834 10260
rect 45554 10248 45560 10260
rect 40828 10220 45560 10248
rect 40828 10208 40834 10220
rect 45554 10208 45560 10220
rect 45612 10208 45618 10260
rect 48038 10208 48044 10260
rect 48096 10248 48102 10260
rect 48317 10251 48375 10257
rect 48317 10248 48329 10251
rect 48096 10220 48329 10248
rect 48096 10208 48102 10220
rect 48317 10217 48329 10220
rect 48363 10217 48375 10251
rect 48317 10211 48375 10217
rect 52365 10251 52423 10257
rect 52365 10217 52377 10251
rect 52411 10217 52423 10251
rect 52365 10211 52423 10217
rect 52825 10251 52883 10257
rect 52825 10217 52837 10251
rect 52871 10248 52883 10251
rect 53926 10248 53932 10260
rect 52871 10220 53932 10248
rect 52871 10217 52883 10220
rect 52825 10211 52883 10217
rect 33229 10183 33287 10189
rect 33229 10180 33241 10183
rect 32416 10152 33241 10180
rect 33229 10149 33241 10152
rect 33275 10180 33287 10183
rect 33318 10180 33324 10192
rect 33275 10152 33324 10180
rect 33275 10149 33287 10152
rect 33229 10143 33287 10149
rect 33318 10140 33324 10152
rect 33376 10140 33382 10192
rect 41414 10180 41420 10192
rect 38672 10152 41420 10180
rect 38672 10124 38700 10152
rect 41414 10140 41420 10152
rect 41472 10140 41478 10192
rect 31481 10115 31539 10121
rect 31481 10081 31493 10115
rect 31527 10081 31539 10115
rect 31481 10075 31539 10081
rect 31846 10072 31852 10124
rect 31904 10112 31910 10124
rect 31904 10084 32996 10112
rect 31904 10072 31910 10084
rect 21082 10004 21088 10056
rect 21140 10044 21146 10056
rect 21177 10047 21235 10053
rect 21177 10044 21189 10047
rect 21140 10016 21189 10044
rect 21140 10004 21146 10016
rect 21177 10013 21189 10016
rect 21223 10013 21235 10047
rect 21177 10007 21235 10013
rect 22094 10004 22100 10056
rect 22152 10044 22158 10056
rect 22152 10016 22197 10044
rect 22152 10004 22158 10016
rect 20456 9948 22094 9976
rect 20349 9939 20407 9945
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 15565 9911 15623 9917
rect 15565 9908 15577 9911
rect 13872 9880 15577 9908
rect 13872 9868 13878 9880
rect 15565 9877 15577 9880
rect 15611 9908 15623 9911
rect 15746 9908 15752 9920
rect 15611 9880 15752 9908
rect 15611 9877 15623 9880
rect 15565 9871 15623 9877
rect 15746 9868 15752 9880
rect 15804 9908 15810 9920
rect 17497 9911 17555 9917
rect 17497 9908 17509 9911
rect 15804 9880 17509 9908
rect 15804 9868 15810 9880
rect 17497 9877 17509 9880
rect 17543 9908 17555 9911
rect 18598 9908 18604 9920
rect 17543 9880 18604 9908
rect 17543 9877 17555 9880
rect 17497 9871 17555 9877
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 18693 9911 18751 9917
rect 18693 9877 18705 9911
rect 18739 9908 18751 9911
rect 18782 9908 18788 9920
rect 18739 9880 18788 9908
rect 18739 9877 18751 9880
rect 18693 9871 18751 9877
rect 18782 9868 18788 9880
rect 18840 9868 18846 9920
rect 20254 9908 20260 9920
rect 20215 9880 20260 9908
rect 20254 9868 20260 9880
rect 20312 9868 20318 9920
rect 22066 9908 22094 9948
rect 24670 9936 24676 9988
rect 24728 9976 24734 9988
rect 24857 9979 24915 9985
rect 24857 9976 24869 9979
rect 24728 9948 24869 9976
rect 24728 9936 24734 9948
rect 24857 9945 24869 9948
rect 24903 9976 24915 9979
rect 27172 9976 27200 10072
rect 30466 10044 30472 10056
rect 30427 10016 30472 10044
rect 30466 10004 30472 10016
rect 30524 10004 30530 10056
rect 31396 10047 31454 10053
rect 31396 10013 31408 10047
rect 31442 10038 31454 10047
rect 31754 10044 31760 10056
rect 31588 10038 31760 10044
rect 31442 10016 31760 10038
rect 31442 10013 31616 10016
rect 31396 10010 31616 10013
rect 31396 10007 31454 10010
rect 31754 10004 31760 10016
rect 31812 10044 31818 10056
rect 32677 10047 32735 10053
rect 32677 10044 32689 10047
rect 31812 10016 32689 10044
rect 31812 10004 31818 10016
rect 32677 10013 32689 10016
rect 32723 10013 32735 10047
rect 32968 10044 32996 10084
rect 33686 10072 33692 10124
rect 33744 10112 33750 10124
rect 34698 10112 34704 10124
rect 33744 10084 34704 10112
rect 33744 10072 33750 10084
rect 34698 10072 34704 10084
rect 34756 10112 34762 10124
rect 35066 10112 35072 10124
rect 34756 10084 35072 10112
rect 34756 10072 34762 10084
rect 35066 10072 35072 10084
rect 35124 10072 35130 10124
rect 36906 10112 36912 10124
rect 36867 10084 36912 10112
rect 36906 10072 36912 10084
rect 36964 10072 36970 10124
rect 38654 10112 38660 10124
rect 38615 10084 38660 10112
rect 38654 10072 38660 10084
rect 38712 10072 38718 10124
rect 40034 10112 40040 10124
rect 39995 10084 40040 10112
rect 40034 10072 40040 10084
rect 40092 10072 40098 10124
rect 40218 10072 40224 10124
rect 40276 10112 40282 10124
rect 41230 10112 41236 10124
rect 40276 10084 41236 10112
rect 40276 10072 40282 10084
rect 41230 10072 41236 10084
rect 41288 10112 41294 10124
rect 43257 10115 43315 10121
rect 43257 10112 43269 10115
rect 41288 10084 43269 10112
rect 41288 10072 41294 10084
rect 43257 10081 43269 10084
rect 43303 10081 43315 10115
rect 51074 10112 51080 10124
rect 50987 10084 51080 10112
rect 43257 10075 43315 10081
rect 51074 10072 51080 10084
rect 51132 10112 51138 10124
rect 52380 10112 52408 10211
rect 53926 10208 53932 10220
rect 53984 10208 53990 10260
rect 55398 10140 55404 10192
rect 55456 10180 55462 10192
rect 55861 10183 55919 10189
rect 55861 10180 55873 10183
rect 55456 10152 55873 10180
rect 55456 10140 55462 10152
rect 55861 10149 55873 10152
rect 55907 10180 55919 10183
rect 55907 10152 56732 10180
rect 55907 10149 55919 10152
rect 55861 10143 55919 10149
rect 51132 10084 52408 10112
rect 52457 10115 52515 10121
rect 51132 10072 51138 10084
rect 52457 10081 52469 10115
rect 52503 10081 52515 10115
rect 55122 10112 55128 10124
rect 52457 10075 52515 10081
rect 52656 10084 55128 10112
rect 39114 10044 39120 10056
rect 32968 10016 34744 10044
rect 39075 10016 39120 10044
rect 32677 10007 32735 10013
rect 24903 9948 27200 9976
rect 24903 9945 24915 9948
rect 24857 9939 24915 9945
rect 28718 9936 28724 9988
rect 28776 9976 28782 9988
rect 29549 9979 29607 9985
rect 29549 9976 29561 9979
rect 28776 9948 29561 9976
rect 28776 9936 28782 9948
rect 29549 9945 29561 9948
rect 29595 9945 29607 9979
rect 31662 9976 31668 9988
rect 31623 9948 31668 9976
rect 29549 9939 29607 9945
rect 31662 9936 31668 9948
rect 31720 9936 31726 9988
rect 32217 9979 32275 9985
rect 32217 9945 32229 9979
rect 32263 9976 32275 9979
rect 33134 9976 33140 9988
rect 32263 9948 33140 9976
rect 32263 9945 32275 9948
rect 32217 9939 32275 9945
rect 26418 9908 26424 9920
rect 22066 9880 26424 9908
rect 26418 9868 26424 9880
rect 26476 9868 26482 9920
rect 30834 9868 30840 9920
rect 30892 9908 30898 9920
rect 32232 9908 32260 9939
rect 33134 9936 33140 9948
rect 33192 9936 33198 9988
rect 34057 9979 34115 9985
rect 34057 9945 34069 9979
rect 34103 9976 34115 9979
rect 34606 9976 34612 9988
rect 34103 9948 34612 9976
rect 34103 9945 34115 9948
rect 34057 9939 34115 9945
rect 34606 9936 34612 9948
rect 34664 9936 34670 9988
rect 30892 9880 32260 9908
rect 33965 9911 34023 9917
rect 30892 9868 30898 9880
rect 33965 9877 33977 9911
rect 34011 9908 34023 9911
rect 34330 9908 34336 9920
rect 34011 9880 34336 9908
rect 34011 9877 34023 9880
rect 33965 9871 34023 9877
rect 34330 9868 34336 9880
rect 34388 9868 34394 9920
rect 34716 9908 34744 10016
rect 39114 10004 39120 10016
rect 39172 10004 39178 10056
rect 39298 10044 39304 10056
rect 39259 10016 39304 10044
rect 39298 10004 39304 10016
rect 39356 10004 39362 10056
rect 51350 10044 51356 10056
rect 51311 10016 51356 10044
rect 51350 10004 51356 10016
rect 51408 10004 51414 10056
rect 52362 10044 52368 10056
rect 52323 10016 52368 10044
rect 52362 10004 52368 10016
rect 52420 10004 52426 10056
rect 36262 9976 36268 9988
rect 36202 9948 36268 9976
rect 36262 9936 36268 9948
rect 36320 9936 36326 9988
rect 37185 9979 37243 9985
rect 37185 9945 37197 9979
rect 37231 9945 37243 9979
rect 37185 9939 37243 9945
rect 36449 9911 36507 9917
rect 36449 9908 36461 9911
rect 34716 9880 36461 9908
rect 36449 9877 36461 9880
rect 36495 9877 36507 9911
rect 37200 9908 37228 9939
rect 38194 9936 38200 9988
rect 38252 9936 38258 9988
rect 38470 9936 38476 9988
rect 38528 9976 38534 9988
rect 39209 9979 39267 9985
rect 39209 9976 39221 9979
rect 38528 9948 39221 9976
rect 38528 9936 38534 9948
rect 39209 9945 39221 9948
rect 39255 9945 39267 9979
rect 39209 9939 39267 9945
rect 42518 9936 42524 9988
rect 42576 9936 42582 9988
rect 42702 9936 42708 9988
rect 42760 9976 42766 9988
rect 42981 9979 43039 9985
rect 42981 9976 42993 9979
rect 42760 9948 42993 9976
rect 42760 9936 42766 9948
rect 42981 9945 42993 9948
rect 43027 9945 43039 9979
rect 45462 9976 45468 9988
rect 45423 9948 45468 9976
rect 42981 9939 43039 9945
rect 45462 9936 45468 9948
rect 45520 9936 45526 9988
rect 51902 9936 51908 9988
rect 51960 9976 51966 9988
rect 52472 9976 52500 10075
rect 52656 10056 52684 10084
rect 55122 10072 55128 10084
rect 55180 10112 55186 10124
rect 56321 10115 56379 10121
rect 56321 10112 56333 10115
rect 55180 10084 56333 10112
rect 55180 10072 55186 10084
rect 56321 10081 56333 10084
rect 56367 10081 56379 10115
rect 56321 10075 56379 10081
rect 56594 10072 56600 10124
rect 56652 10072 56658 10124
rect 56704 10112 56732 10152
rect 57330 10112 57336 10124
rect 56704 10084 57336 10112
rect 57330 10072 57336 10084
rect 57388 10112 57394 10124
rect 58069 10115 58127 10121
rect 58069 10112 58081 10115
rect 57388 10084 58081 10112
rect 57388 10072 57394 10084
rect 58069 10081 58081 10084
rect 58115 10081 58127 10115
rect 58069 10075 58127 10081
rect 52638 10044 52644 10056
rect 52551 10016 52644 10044
rect 52638 10004 52644 10016
rect 52696 10004 52702 10056
rect 56612 10044 56640 10072
rect 56612 10016 56718 10044
rect 51960 9948 52500 9976
rect 51960 9936 51966 9948
rect 57514 9936 57520 9988
rect 57572 9976 57578 9988
rect 57793 9979 57851 9985
rect 57793 9976 57805 9979
rect 57572 9948 57805 9976
rect 57572 9936 57578 9948
rect 57793 9945 57805 9948
rect 57839 9945 57851 9979
rect 57793 9939 57851 9945
rect 38102 9908 38108 9920
rect 37200 9880 38108 9908
rect 36449 9871 36507 9877
rect 38102 9868 38108 9880
rect 38160 9868 38166 9920
rect 40126 9908 40132 9920
rect 40087 9880 40132 9908
rect 40126 9868 40132 9880
rect 40184 9868 40190 9920
rect 40221 9911 40279 9917
rect 40221 9877 40233 9911
rect 40267 9908 40279 9911
rect 41138 9908 41144 9920
rect 40267 9880 41144 9908
rect 40267 9877 40279 9880
rect 40221 9871 40279 9877
rect 41138 9868 41144 9880
rect 41196 9868 41202 9920
rect 41230 9868 41236 9920
rect 41288 9908 41294 9920
rect 41509 9911 41567 9917
rect 41509 9908 41521 9911
rect 41288 9880 41521 9908
rect 41288 9868 41294 9880
rect 41509 9877 41521 9880
rect 41555 9877 41567 9911
rect 41509 9871 41567 9877
rect 43809 9911 43867 9917
rect 43809 9877 43821 9911
rect 43855 9908 43867 9911
rect 44174 9908 44180 9920
rect 43855 9880 44180 9908
rect 43855 9877 43867 9880
rect 43809 9871 43867 9877
rect 44174 9868 44180 9880
rect 44232 9908 44238 9920
rect 44269 9911 44327 9917
rect 44269 9908 44281 9911
rect 44232 9880 44281 9908
rect 44232 9868 44238 9880
rect 44269 9877 44281 9880
rect 44315 9877 44327 9911
rect 44269 9871 44327 9877
rect 1104 9818 58880 9840
rect 1104 9766 15398 9818
rect 15450 9766 15462 9818
rect 15514 9766 15526 9818
rect 15578 9766 15590 9818
rect 15642 9766 15654 9818
rect 15706 9766 29846 9818
rect 29898 9766 29910 9818
rect 29962 9766 29974 9818
rect 30026 9766 30038 9818
rect 30090 9766 30102 9818
rect 30154 9766 44294 9818
rect 44346 9766 44358 9818
rect 44410 9766 44422 9818
rect 44474 9766 44486 9818
rect 44538 9766 44550 9818
rect 44602 9766 58880 9818
rect 1104 9744 58880 9766
rect 17586 9664 17592 9716
rect 17644 9704 17650 9716
rect 20254 9704 20260 9716
rect 17644 9676 18000 9704
rect 17644 9664 17650 9676
rect 17972 9636 18000 9676
rect 19076 9676 20260 9704
rect 19076 9636 19104 9676
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 20438 9664 20444 9716
rect 20496 9704 20502 9716
rect 21910 9704 21916 9716
rect 20496 9676 21916 9704
rect 20496 9664 20502 9676
rect 21910 9664 21916 9676
rect 21968 9704 21974 9716
rect 30650 9704 30656 9716
rect 21968 9676 22061 9704
rect 27448 9676 30656 9704
rect 21968 9664 21974 9676
rect 20714 9636 20720 9648
rect 17972 9608 19182 9636
rect 20675 9608 20720 9636
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 21821 9639 21879 9645
rect 21821 9605 21833 9639
rect 21867 9636 21879 9639
rect 21928 9636 21956 9664
rect 21867 9608 21956 9636
rect 21867 9605 21879 9608
rect 21821 9599 21879 9605
rect 22462 9596 22468 9648
rect 22520 9636 22526 9648
rect 25869 9639 25927 9645
rect 25869 9636 25881 9639
rect 22520 9608 25881 9636
rect 22520 9596 22526 9608
rect 25869 9605 25881 9608
rect 25915 9605 25927 9639
rect 25869 9599 25927 9605
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9568 20867 9571
rect 23842 9568 23848 9580
rect 20855 9540 23848 9568
rect 20855 9537 20867 9540
rect 20809 9531 20867 9537
rect 23842 9528 23848 9540
rect 23900 9528 23906 9580
rect 18414 9500 18420 9512
rect 17880 9472 18420 9500
rect 17770 9432 17776 9444
rect 12406 9404 17776 9432
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 12406 9364 12434 9404
rect 17770 9392 17776 9404
rect 17828 9392 17834 9444
rect 3292 9336 12434 9364
rect 3292 9324 3298 9336
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 17880 9373 17908 9472
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 18690 9500 18696 9512
rect 18651 9472 18696 9500
rect 18690 9460 18696 9472
rect 18748 9460 18754 9512
rect 24670 9500 24676 9512
rect 24631 9472 24676 9500
rect 24670 9460 24676 9472
rect 24728 9460 24734 9512
rect 27448 9509 27476 9676
rect 30650 9664 30656 9676
rect 30708 9664 30714 9716
rect 34606 9664 34612 9716
rect 34664 9704 34670 9716
rect 36262 9704 36268 9716
rect 34664 9676 36268 9704
rect 34664 9664 34670 9676
rect 28442 9596 28448 9648
rect 28500 9636 28506 9648
rect 28629 9639 28687 9645
rect 28629 9636 28641 9639
rect 28500 9608 28641 9636
rect 28500 9596 28506 9608
rect 28629 9605 28641 9608
rect 28675 9605 28687 9639
rect 28629 9599 28687 9605
rect 29270 9596 29276 9648
rect 29328 9636 29334 9648
rect 29917 9639 29975 9645
rect 29917 9636 29929 9639
rect 29328 9608 29929 9636
rect 29328 9596 29334 9608
rect 29917 9605 29929 9608
rect 29963 9605 29975 9639
rect 35268 9636 35296 9676
rect 36262 9664 36268 9676
rect 36320 9664 36326 9716
rect 40126 9664 40132 9716
rect 40184 9704 40190 9716
rect 40747 9707 40805 9713
rect 40747 9704 40759 9707
rect 40184 9676 40759 9704
rect 40184 9664 40190 9676
rect 40747 9673 40759 9676
rect 40793 9704 40805 9707
rect 42610 9704 42616 9716
rect 40793 9676 42616 9704
rect 40793 9673 40805 9676
rect 40747 9667 40805 9673
rect 42610 9664 42616 9676
rect 42668 9664 42674 9716
rect 43530 9704 43536 9716
rect 43491 9676 43536 9704
rect 43530 9664 43536 9676
rect 43588 9664 43594 9716
rect 49786 9704 49792 9716
rect 49528 9676 49792 9704
rect 38378 9636 38384 9648
rect 35190 9608 35296 9636
rect 38339 9608 38384 9636
rect 29917 9599 29975 9605
rect 38378 9596 38384 9608
rect 38436 9596 38442 9648
rect 40034 9596 40040 9648
rect 40092 9636 40098 9648
rect 40957 9639 41015 9645
rect 40957 9636 40969 9639
rect 40092 9608 40969 9636
rect 40092 9596 40098 9608
rect 40957 9605 40969 9608
rect 41003 9636 41015 9639
rect 41230 9636 41236 9648
rect 41003 9608 41236 9636
rect 41003 9605 41015 9608
rect 40957 9599 41015 9605
rect 41230 9596 41236 9608
rect 41288 9596 41294 9648
rect 41601 9639 41659 9645
rect 41601 9605 41613 9639
rect 41647 9636 41659 9639
rect 43548 9636 43576 9664
rect 41647 9608 43576 9636
rect 41647 9605 41659 9608
rect 41601 9599 41659 9605
rect 44818 9596 44824 9648
rect 44876 9636 44882 9648
rect 49528 9636 49556 9676
rect 49786 9664 49792 9676
rect 49844 9664 49850 9716
rect 57514 9664 57520 9716
rect 57572 9704 57578 9716
rect 57572 9676 58112 9704
rect 57572 9664 57578 9676
rect 44876 9608 47808 9636
rect 44876 9596 44882 9608
rect 31938 9528 31944 9580
rect 31996 9568 32002 9580
rect 32677 9571 32735 9577
rect 32677 9568 32689 9571
rect 31996 9540 32689 9568
rect 31996 9528 32002 9540
rect 32677 9537 32689 9540
rect 32723 9537 32735 9571
rect 33686 9568 33692 9580
rect 33647 9540 33692 9568
rect 32677 9531 32735 9537
rect 33686 9528 33692 9540
rect 33744 9528 33750 9580
rect 35986 9528 35992 9580
rect 36044 9568 36050 9580
rect 36173 9571 36231 9577
rect 36173 9568 36185 9571
rect 36044 9540 36185 9568
rect 36044 9528 36050 9540
rect 36173 9537 36185 9540
rect 36219 9537 36231 9571
rect 36173 9531 36231 9537
rect 36906 9528 36912 9580
rect 36964 9568 36970 9580
rect 37461 9571 37519 9577
rect 37461 9568 37473 9571
rect 36964 9540 37473 9568
rect 36964 9528 36970 9540
rect 37461 9537 37473 9540
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 41322 9528 41328 9580
rect 41380 9568 41386 9580
rect 42613 9571 42671 9577
rect 42613 9568 42625 9571
rect 41380 9540 42625 9568
rect 41380 9528 41386 9540
rect 42613 9537 42625 9540
rect 42659 9537 42671 9571
rect 42613 9531 42671 9537
rect 44453 9571 44511 9577
rect 44453 9537 44465 9571
rect 44499 9568 44511 9571
rect 44726 9568 44732 9580
rect 44499 9540 44732 9568
rect 44499 9537 44511 9540
rect 44453 9531 44511 9537
rect 44726 9528 44732 9540
rect 44784 9568 44790 9580
rect 45462 9568 45468 9580
rect 44784 9540 45468 9568
rect 44784 9528 44790 9540
rect 45462 9528 45468 9540
rect 45520 9528 45526 9580
rect 47780 9577 47808 9608
rect 48884 9608 49556 9636
rect 47765 9571 47823 9577
rect 47765 9537 47777 9571
rect 47811 9568 47823 9571
rect 48222 9568 48228 9580
rect 47811 9540 48228 9568
rect 47811 9537 47823 9540
rect 47765 9531 47823 9537
rect 48222 9528 48228 9540
rect 48280 9528 48286 9580
rect 48884 9577 48912 9608
rect 51442 9596 51448 9648
rect 51500 9636 51506 9648
rect 51813 9639 51871 9645
rect 51813 9636 51825 9639
rect 51500 9608 51825 9636
rect 51500 9596 51506 9608
rect 51813 9605 51825 9608
rect 51859 9605 51871 9639
rect 51813 9599 51871 9605
rect 51997 9639 52055 9645
rect 51997 9605 52009 9639
rect 52043 9636 52055 9639
rect 52638 9636 52644 9648
rect 52043 9608 52644 9636
rect 52043 9605 52055 9608
rect 51997 9599 52055 9605
rect 52638 9596 52644 9608
rect 52696 9596 52702 9648
rect 54570 9636 54576 9648
rect 54531 9608 54576 9636
rect 54570 9596 54576 9608
rect 54628 9596 54634 9648
rect 56594 9636 56600 9648
rect 55798 9608 56600 9636
rect 56594 9596 56600 9608
rect 56652 9596 56658 9648
rect 58084 9645 58112 9676
rect 58069 9639 58127 9645
rect 58069 9605 58081 9639
rect 58115 9605 58127 9639
rect 58069 9599 58127 9605
rect 48869 9571 48927 9577
rect 48869 9537 48881 9571
rect 48915 9537 48927 9571
rect 48869 9531 48927 9537
rect 50246 9528 50252 9580
rect 50304 9528 50310 9580
rect 54294 9568 54300 9580
rect 54255 9540 54300 9568
rect 54294 9528 54300 9540
rect 54352 9528 54358 9580
rect 26053 9503 26111 9509
rect 26053 9469 26065 9503
rect 26099 9469 26111 9503
rect 26053 9463 26111 9469
rect 27433 9503 27491 9509
rect 27433 9469 27445 9503
rect 27479 9469 27491 9503
rect 27433 9463 27491 9469
rect 26068 9432 26096 9463
rect 28074 9460 28080 9512
rect 28132 9500 28138 9512
rect 28813 9503 28871 9509
rect 28813 9500 28825 9503
rect 28132 9472 28825 9500
rect 28132 9460 28138 9472
rect 28813 9469 28825 9472
rect 28859 9469 28871 9503
rect 28813 9463 28871 9469
rect 29733 9503 29791 9509
rect 29733 9469 29745 9503
rect 29779 9500 29791 9503
rect 30558 9500 30564 9512
rect 29779 9472 30564 9500
rect 29779 9469 29791 9472
rect 29733 9463 29791 9469
rect 30558 9460 30564 9472
rect 30616 9460 30622 9512
rect 30650 9460 30656 9512
rect 30708 9500 30714 9512
rect 33962 9500 33968 9512
rect 30708 9472 30753 9500
rect 33923 9472 33968 9500
rect 30708 9460 30714 9472
rect 33962 9460 33968 9472
rect 34020 9460 34026 9512
rect 37277 9503 37335 9509
rect 37277 9500 37289 9503
rect 35084 9472 37289 9500
rect 35084 9444 35112 9472
rect 37277 9469 37289 9472
rect 37323 9500 37335 9503
rect 38838 9500 38844 9512
rect 37323 9472 38844 9500
rect 37323 9469 37335 9472
rect 37277 9463 37335 9469
rect 38838 9460 38844 9472
rect 38896 9460 38902 9512
rect 40954 9460 40960 9512
rect 41012 9500 41018 9512
rect 42521 9503 42579 9509
rect 42521 9500 42533 9503
rect 41012 9472 42533 9500
rect 41012 9460 41018 9472
rect 42521 9469 42533 9472
rect 42567 9469 42579 9503
rect 42521 9463 42579 9469
rect 47857 9503 47915 9509
rect 47857 9469 47869 9503
rect 47903 9500 47915 9503
rect 48314 9500 48320 9512
rect 47903 9472 48320 9500
rect 47903 9469 47915 9472
rect 47857 9463 47915 9469
rect 48314 9460 48320 9472
rect 48372 9460 48378 9512
rect 49145 9503 49203 9509
rect 49145 9500 49157 9503
rect 48976 9472 49157 9500
rect 27982 9432 27988 9444
rect 26068 9404 27988 9432
rect 27982 9392 27988 9404
rect 28040 9392 28046 9444
rect 31754 9392 31760 9444
rect 31812 9432 31818 9444
rect 32493 9435 32551 9441
rect 32493 9432 32505 9435
rect 31812 9404 32505 9432
rect 31812 9392 31818 9404
rect 32493 9401 32505 9404
rect 32539 9401 32551 9435
rect 33686 9432 33692 9444
rect 32493 9395 32551 9401
rect 33244 9404 33692 9432
rect 17865 9367 17923 9373
rect 17865 9364 17877 9367
rect 16356 9336 17877 9364
rect 16356 9324 16362 9336
rect 17865 9333 17877 9336
rect 17911 9333 17923 9367
rect 17865 9327 17923 9333
rect 20165 9367 20223 9373
rect 20165 9333 20177 9367
rect 20211 9364 20223 9367
rect 20254 9364 20260 9376
rect 20211 9336 20260 9364
rect 20211 9333 20223 9336
rect 20165 9327 20223 9333
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 27246 9324 27252 9376
rect 27304 9364 27310 9376
rect 28166 9364 28172 9376
rect 27304 9336 28172 9364
rect 27304 9324 27310 9336
rect 28166 9324 28172 9336
rect 28224 9364 28230 9376
rect 30190 9364 30196 9376
rect 28224 9336 30196 9364
rect 28224 9324 28230 9336
rect 30190 9324 30196 9336
rect 30248 9324 30254 9376
rect 30374 9324 30380 9376
rect 30432 9364 30438 9376
rect 33244 9364 33272 9404
rect 33686 9392 33692 9404
rect 33744 9392 33750 9444
rect 35066 9392 35072 9444
rect 35124 9392 35130 9444
rect 35894 9392 35900 9444
rect 35952 9432 35958 9444
rect 35989 9435 36047 9441
rect 35989 9432 36001 9435
rect 35952 9404 36001 9432
rect 35952 9392 35958 9404
rect 35989 9401 36001 9404
rect 36035 9401 36047 9435
rect 35989 9395 36047 9401
rect 39298 9392 39304 9444
rect 39356 9432 39362 9444
rect 40589 9435 40647 9441
rect 40589 9432 40601 9435
rect 39356 9404 40601 9432
rect 39356 9392 39362 9404
rect 40589 9401 40601 9404
rect 40635 9401 40647 9435
rect 44637 9435 44695 9441
rect 44637 9432 44649 9435
rect 40589 9395 40647 9401
rect 40696 9404 44649 9432
rect 30432 9336 33272 9364
rect 30432 9324 30438 9336
rect 33318 9324 33324 9376
rect 33376 9364 33382 9376
rect 35437 9367 35495 9373
rect 35437 9364 35449 9367
rect 33376 9336 35449 9364
rect 33376 9324 33382 9336
rect 35437 9333 35449 9336
rect 35483 9333 35495 9367
rect 35437 9327 35495 9333
rect 38930 9324 38936 9376
rect 38988 9364 38994 9376
rect 39669 9367 39727 9373
rect 39669 9364 39681 9367
rect 38988 9336 39681 9364
rect 38988 9324 38994 9336
rect 39669 9333 39681 9336
rect 39715 9333 39727 9367
rect 39669 9327 39727 9333
rect 39758 9324 39764 9376
rect 39816 9364 39822 9376
rect 40696 9364 40724 9404
rect 44637 9401 44649 9404
rect 44683 9432 44695 9435
rect 46934 9432 46940 9444
rect 44683 9404 46940 9432
rect 44683 9401 44695 9404
rect 44637 9395 44695 9401
rect 46934 9392 46940 9404
rect 46992 9392 46998 9444
rect 48133 9435 48191 9441
rect 48133 9401 48145 9435
rect 48179 9432 48191 9435
rect 48976 9432 49004 9472
rect 49145 9469 49157 9472
rect 49191 9469 49203 9503
rect 49145 9463 49203 9469
rect 50617 9503 50675 9509
rect 50617 9469 50629 9503
rect 50663 9500 50675 9503
rect 51074 9500 51080 9512
rect 50663 9472 51080 9500
rect 50663 9469 50675 9472
rect 50617 9463 50675 9469
rect 51074 9460 51080 9472
rect 51132 9460 51138 9512
rect 56042 9500 56048 9512
rect 56003 9472 56048 9500
rect 56042 9460 56048 9472
rect 56100 9460 56106 9512
rect 48179 9404 49004 9432
rect 48179 9401 48191 9404
rect 48133 9395 48191 9401
rect 39816 9336 40724 9364
rect 40773 9367 40831 9373
rect 39816 9324 39822 9336
rect 40773 9333 40785 9367
rect 40819 9364 40831 9367
rect 40862 9364 40868 9376
rect 40819 9336 40868 9364
rect 40819 9333 40831 9336
rect 40773 9327 40831 9333
rect 40862 9324 40868 9336
rect 40920 9324 40926 9376
rect 41046 9324 41052 9376
rect 41104 9364 41110 9376
rect 41509 9367 41567 9373
rect 41509 9364 41521 9367
rect 41104 9336 41521 9364
rect 41104 9324 41110 9336
rect 41509 9333 41521 9336
rect 41555 9333 41567 9367
rect 42886 9364 42892 9376
rect 42847 9336 42892 9364
rect 41509 9327 41567 9333
rect 42886 9324 42892 9336
rect 42944 9324 42950 9376
rect 1104 9274 58880 9296
rect 1104 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 8302 9274
rect 8354 9222 8366 9274
rect 8418 9222 8430 9274
rect 8482 9222 22622 9274
rect 22674 9222 22686 9274
rect 22738 9222 22750 9274
rect 22802 9222 22814 9274
rect 22866 9222 22878 9274
rect 22930 9222 37070 9274
rect 37122 9222 37134 9274
rect 37186 9222 37198 9274
rect 37250 9222 37262 9274
rect 37314 9222 37326 9274
rect 37378 9222 51518 9274
rect 51570 9222 51582 9274
rect 51634 9222 51646 9274
rect 51698 9222 51710 9274
rect 51762 9222 51774 9274
rect 51826 9222 58880 9274
rect 1104 9200 58880 9222
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 18601 9163 18659 9169
rect 18601 9129 18613 9163
rect 18647 9160 18659 9163
rect 18690 9160 18696 9172
rect 18647 9132 18696 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 19521 9163 19579 9169
rect 19521 9129 19533 9163
rect 19567 9160 19579 9163
rect 19886 9160 19892 9172
rect 19567 9132 19892 9160
rect 19567 9129 19579 9132
rect 19521 9123 19579 9129
rect 19886 9120 19892 9132
rect 19944 9120 19950 9172
rect 20990 9160 20996 9172
rect 20951 9132 20996 9160
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 26697 9163 26755 9169
rect 26697 9129 26709 9163
rect 26743 9160 26755 9163
rect 33962 9160 33968 9172
rect 26743 9132 33968 9160
rect 26743 9129 26755 9132
rect 26697 9123 26755 9129
rect 33962 9120 33968 9132
rect 34020 9120 34026 9172
rect 34146 9120 34152 9172
rect 34204 9160 34210 9172
rect 35161 9163 35219 9169
rect 35161 9160 35173 9163
rect 34204 9132 35173 9160
rect 34204 9120 34210 9132
rect 35161 9129 35173 9132
rect 35207 9129 35219 9163
rect 38562 9160 38568 9172
rect 35161 9123 35219 9129
rect 36096 9132 38568 9160
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 3252 8956 3280 9120
rect 20254 9092 20260 9104
rect 20215 9064 20260 9092
rect 20254 9052 20260 9064
rect 20312 9052 20318 9104
rect 25777 9095 25835 9101
rect 25777 9061 25789 9095
rect 25823 9092 25835 9095
rect 27246 9092 27252 9104
rect 25823 9064 27252 9092
rect 25823 9061 25835 9064
rect 25777 9055 25835 9061
rect 27246 9052 27252 9064
rect 27304 9052 27310 9104
rect 30101 9095 30159 9101
rect 28276 9064 30052 9092
rect 28276 9033 28304 9064
rect 26513 9027 26571 9033
rect 26513 8993 26525 9027
rect 26559 9024 26571 9027
rect 27341 9027 27399 9033
rect 27341 9024 27353 9027
rect 26559 8996 27353 9024
rect 26559 8993 26571 8996
rect 26513 8987 26571 8993
rect 27341 8993 27353 8996
rect 27387 8993 27399 9027
rect 27341 8987 27399 8993
rect 27893 9027 27951 9033
rect 27893 8993 27905 9027
rect 27939 8993 27951 9027
rect 27893 8987 27951 8993
rect 28261 9027 28319 9033
rect 28261 8993 28273 9027
rect 28307 8993 28319 9027
rect 28261 8987 28319 8993
rect 28353 9027 28411 9033
rect 28353 8993 28365 9027
rect 28399 9024 28411 9027
rect 29362 9024 29368 9036
rect 28399 8996 29368 9024
rect 28399 8993 28411 8996
rect 28353 8987 28411 8993
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 2731 8928 3280 8956
rect 16316 8928 16865 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 16316 8832 16344 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 26418 8956 26424 8968
rect 26379 8928 26424 8956
rect 16853 8919 16911 8925
rect 26418 8916 26424 8928
rect 26476 8916 26482 8968
rect 27246 8956 27252 8968
rect 27207 8928 27252 8956
rect 27246 8916 27252 8928
rect 27304 8916 27310 8968
rect 27433 8959 27491 8965
rect 27433 8925 27445 8959
rect 27479 8956 27491 8959
rect 27908 8956 27936 8987
rect 29362 8984 29368 8996
rect 29420 8984 29426 9036
rect 29638 9024 29644 9036
rect 29599 8996 29644 9024
rect 29638 8984 29644 8996
rect 29696 8984 29702 9036
rect 28077 8959 28135 8965
rect 28077 8956 28089 8959
rect 27479 8928 27936 8956
rect 28000 8928 28089 8956
rect 27479 8925 27491 8928
rect 27433 8919 27491 8925
rect 17126 8888 17132 8900
rect 17087 8860 17132 8888
rect 17126 8848 17132 8860
rect 17184 8848 17190 8900
rect 17586 8848 17592 8900
rect 17644 8848 17650 8900
rect 19978 8888 19984 8900
rect 19939 8860 19984 8888
rect 19978 8848 19984 8860
rect 20036 8848 20042 8900
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 1728 8792 2513 8820
rect 1728 8780 1734 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 16298 8820 16304 8832
rect 16259 8792 16304 8820
rect 2501 8783 2559 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 20438 8820 20444 8832
rect 20399 8792 20444 8820
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 21174 8780 21180 8832
rect 21232 8820 21238 8832
rect 21453 8823 21511 8829
rect 21453 8820 21465 8823
rect 21232 8792 21465 8820
rect 21232 8780 21238 8792
rect 21453 8789 21465 8792
rect 21499 8789 21511 8823
rect 28000 8820 28028 8928
rect 28077 8925 28089 8928
rect 28123 8925 28135 8959
rect 28077 8919 28135 8925
rect 28166 8916 28172 8968
rect 28224 8956 28230 8968
rect 29730 8956 29736 8968
rect 28224 8928 28269 8956
rect 29691 8928 29736 8956
rect 28224 8916 28230 8928
rect 29730 8916 29736 8928
rect 29788 8916 29794 8968
rect 30024 8956 30052 9064
rect 30101 9061 30113 9095
rect 30147 9092 30159 9095
rect 30147 9064 31754 9092
rect 30147 9061 30159 9064
rect 30101 9055 30159 9061
rect 30466 8984 30472 9036
rect 30524 9024 30530 9036
rect 31021 9027 31079 9033
rect 31021 9024 31033 9027
rect 30524 8996 31033 9024
rect 30524 8984 30530 8996
rect 31021 8993 31033 8996
rect 31067 8993 31079 9027
rect 31570 9024 31576 9036
rect 31021 8987 31079 8993
rect 31128 8996 31576 9024
rect 31128 8956 31156 8996
rect 31570 8984 31576 8996
rect 31628 8984 31634 9036
rect 31726 9024 31754 9064
rect 33686 9052 33692 9104
rect 33744 9092 33750 9104
rect 35066 9092 35072 9104
rect 33744 9064 35072 9092
rect 33744 9052 33750 9064
rect 35066 9052 35072 9064
rect 35124 9052 35130 9104
rect 34882 9024 34888 9036
rect 31726 8996 34888 9024
rect 34882 8984 34888 8996
rect 34940 8984 34946 9036
rect 30024 8928 31156 8956
rect 31389 8959 31447 8965
rect 31389 8925 31401 8959
rect 31435 8956 31447 8959
rect 31938 8956 31944 8968
rect 31435 8928 31944 8956
rect 31435 8925 31447 8928
rect 31389 8919 31447 8925
rect 31938 8916 31944 8928
rect 31996 8916 32002 8968
rect 32398 8956 32404 8968
rect 32359 8928 32404 8956
rect 32398 8916 32404 8928
rect 32456 8916 32462 8968
rect 35084 8956 35112 9052
rect 35176 9024 35204 9123
rect 36096 9024 36124 9132
rect 38562 9120 38568 9132
rect 38620 9120 38626 9172
rect 40313 9163 40371 9169
rect 40313 9129 40325 9163
rect 40359 9160 40371 9163
rect 40862 9160 40868 9172
rect 40359 9132 40868 9160
rect 40359 9129 40371 9132
rect 40313 9123 40371 9129
rect 40862 9120 40868 9132
rect 40920 9120 40926 9172
rect 41233 9163 41291 9169
rect 41233 9129 41245 9163
rect 41279 9160 41291 9163
rect 41322 9160 41328 9172
rect 41279 9132 41328 9160
rect 41279 9129 41291 9132
rect 41233 9123 41291 9129
rect 36817 9095 36875 9101
rect 36817 9061 36829 9095
rect 36863 9092 36875 9095
rect 38654 9092 38660 9104
rect 36863 9064 38660 9092
rect 36863 9061 36875 9064
rect 36817 9055 36875 9061
rect 38654 9052 38660 9064
rect 38712 9052 38718 9104
rect 38746 9052 38752 9104
rect 38804 9092 38810 9104
rect 38804 9064 38976 9092
rect 38804 9052 38810 9064
rect 35176 8996 36124 9024
rect 35161 8959 35219 8965
rect 35161 8956 35173 8959
rect 35084 8928 35173 8956
rect 35161 8925 35173 8928
rect 35207 8925 35219 8959
rect 35161 8919 35219 8925
rect 35253 8959 35311 8965
rect 35253 8925 35265 8959
rect 35299 8925 35311 8959
rect 35253 8919 35311 8925
rect 28718 8848 28724 8900
rect 28776 8888 28782 8900
rect 28997 8891 29055 8897
rect 28997 8888 29009 8891
rect 28776 8860 29009 8888
rect 28776 8848 28782 8860
rect 28997 8857 29009 8860
rect 29043 8888 29055 8891
rect 31297 8891 31355 8897
rect 31297 8888 31309 8891
rect 29043 8860 31309 8888
rect 29043 8857 29055 8860
rect 28997 8851 29055 8857
rect 31297 8857 31309 8860
rect 31343 8888 31355 8891
rect 31478 8888 31484 8900
rect 31343 8860 31484 8888
rect 31343 8857 31355 8860
rect 31297 8851 31355 8857
rect 31478 8848 31484 8860
rect 31536 8848 31542 8900
rect 32674 8888 32680 8900
rect 32635 8860 32680 8888
rect 32674 8848 32680 8860
rect 32732 8848 32738 8900
rect 34330 8888 34336 8900
rect 33902 8860 34336 8888
rect 34330 8848 34336 8860
rect 34388 8848 34394 8900
rect 34422 8848 34428 8900
rect 34480 8888 34486 8900
rect 35268 8888 35296 8919
rect 35434 8888 35440 8900
rect 34480 8860 35296 8888
rect 35395 8860 35440 8888
rect 34480 8848 34486 8860
rect 35434 8848 35440 8860
rect 35492 8848 35498 8900
rect 36096 8888 36124 8996
rect 38105 9027 38163 9033
rect 38105 8993 38117 9027
rect 38151 9024 38163 9027
rect 38194 9024 38200 9036
rect 38151 8996 38200 9024
rect 38151 8993 38163 8996
rect 38105 8987 38163 8993
rect 38194 8984 38200 8996
rect 38252 8984 38258 9036
rect 38948 9033 38976 9064
rect 38933 9027 38991 9033
rect 38933 8993 38945 9027
rect 38979 9024 38991 9027
rect 39114 9024 39120 9036
rect 38979 8996 39120 9024
rect 38979 8993 38991 8996
rect 38933 8987 38991 8993
rect 39114 8984 39120 8996
rect 39172 9024 39178 9036
rect 40221 9027 40279 9033
rect 40221 9024 40233 9027
rect 39172 8996 40233 9024
rect 39172 8984 39178 8996
rect 40221 8993 40233 8996
rect 40267 9024 40279 9027
rect 41248 9024 41276 9123
rect 41322 9120 41328 9132
rect 41380 9120 41386 9172
rect 42723 9163 42781 9169
rect 42723 9129 42735 9163
rect 42769 9160 42781 9163
rect 42886 9160 42892 9172
rect 42769 9132 42892 9160
rect 42769 9129 42781 9132
rect 42723 9123 42781 9129
rect 42886 9120 42892 9132
rect 42944 9120 42950 9172
rect 48222 9160 48228 9172
rect 48183 9132 48228 9160
rect 48222 9120 48228 9132
rect 48280 9160 48286 9172
rect 50341 9163 50399 9169
rect 50341 9160 50353 9163
rect 48280 9132 50353 9160
rect 48280 9120 48286 9132
rect 50341 9129 50353 9132
rect 50387 9160 50399 9163
rect 50982 9160 50988 9172
rect 50387 9132 50988 9160
rect 50387 9129 50399 9132
rect 50341 9123 50399 9129
rect 50982 9120 50988 9132
rect 51040 9120 51046 9172
rect 55122 9120 55128 9172
rect 55180 9160 55186 9172
rect 55180 9132 56088 9160
rect 55180 9120 55186 9132
rect 43717 9095 43775 9101
rect 43717 9061 43729 9095
rect 43763 9092 43775 9095
rect 45554 9092 45560 9104
rect 43763 9064 45560 9092
rect 43763 9061 43775 9064
rect 43717 9055 43775 9061
rect 45554 9052 45560 9064
rect 45612 9052 45618 9104
rect 40267 8996 41276 9024
rect 40267 8993 40279 8996
rect 40221 8987 40279 8993
rect 42334 8984 42340 9036
rect 42392 9024 42398 9036
rect 42981 9027 43039 9033
rect 42981 9024 42993 9027
rect 42392 8996 42993 9024
rect 42392 8984 42398 8996
rect 42981 8993 42993 8996
rect 43027 8993 43039 9027
rect 42981 8987 43039 8993
rect 45649 9027 45707 9033
rect 45649 8993 45661 9027
rect 45695 9024 45707 9027
rect 46198 9024 46204 9036
rect 45695 8996 46204 9024
rect 45695 8993 45707 8996
rect 45649 8987 45707 8993
rect 46198 8984 46204 8996
rect 46256 8984 46262 9036
rect 56060 9024 56088 9132
rect 57057 9027 57115 9033
rect 57057 9024 57069 9027
rect 56060 8996 57069 9024
rect 57057 8993 57069 8996
rect 57103 8993 57115 9027
rect 57330 9024 57336 9036
rect 57291 8996 57336 9024
rect 57057 8987 57115 8993
rect 57330 8984 57336 8996
rect 57388 8984 57394 9036
rect 36449 8959 36507 8965
rect 36449 8925 36461 8959
rect 36495 8956 36507 8959
rect 37829 8959 37887 8965
rect 36495 8928 37780 8956
rect 36495 8925 36507 8928
rect 36449 8919 36507 8925
rect 36541 8891 36599 8897
rect 36541 8888 36553 8891
rect 36096 8860 36553 8888
rect 36541 8857 36553 8860
rect 36587 8857 36599 8891
rect 37752 8888 37780 8928
rect 37829 8925 37841 8959
rect 37875 8956 37887 8959
rect 38010 8956 38016 8968
rect 37875 8928 38016 8956
rect 37875 8925 37887 8928
rect 37829 8919 37887 8925
rect 38010 8916 38016 8928
rect 38068 8916 38074 8968
rect 38286 8916 38292 8968
rect 38344 8956 38350 8968
rect 38654 8956 38660 8968
rect 38344 8928 38660 8956
rect 38344 8916 38350 8928
rect 38654 8916 38660 8928
rect 38712 8916 38718 8968
rect 38749 8959 38807 8965
rect 38749 8925 38761 8959
rect 38795 8925 38807 8959
rect 38749 8919 38807 8925
rect 38764 8888 38792 8919
rect 38838 8916 38844 8968
rect 38896 8956 38902 8968
rect 39022 8956 39028 8968
rect 38896 8928 38941 8956
rect 38983 8928 39028 8956
rect 38896 8916 38902 8928
rect 39022 8916 39028 8928
rect 39080 8916 39086 8968
rect 40034 8956 40040 8968
rect 39995 8928 40040 8956
rect 40034 8916 40040 8928
rect 40092 8916 40098 8968
rect 40310 8956 40316 8968
rect 40271 8928 40316 8956
rect 40310 8916 40316 8928
rect 40368 8916 40374 8968
rect 43533 8959 43591 8965
rect 43533 8925 43545 8959
rect 43579 8956 43591 8959
rect 44082 8956 44088 8968
rect 43579 8928 44088 8956
rect 43579 8925 43591 8928
rect 43533 8919 43591 8925
rect 44082 8916 44088 8928
rect 44140 8916 44146 8968
rect 45094 8916 45100 8968
rect 45152 8956 45158 8968
rect 45557 8959 45615 8965
rect 45557 8956 45569 8959
rect 45152 8928 45569 8956
rect 45152 8916 45158 8928
rect 45557 8925 45569 8928
rect 45603 8925 45615 8959
rect 45557 8919 45615 8925
rect 50157 8959 50215 8965
rect 50157 8925 50169 8959
rect 50203 8925 50215 8959
rect 50157 8919 50215 8925
rect 39298 8888 39304 8900
rect 37752 8860 39304 8888
rect 36541 8851 36599 8857
rect 39298 8848 39304 8860
rect 39356 8848 39362 8900
rect 42426 8888 42432 8900
rect 42274 8860 42432 8888
rect 42426 8848 42432 8860
rect 42484 8848 42490 8900
rect 44174 8848 44180 8900
rect 44232 8888 44238 8900
rect 44361 8891 44419 8897
rect 44361 8888 44373 8891
rect 44232 8860 44373 8888
rect 44232 8848 44238 8860
rect 44361 8857 44373 8860
rect 44407 8857 44419 8891
rect 45922 8888 45928 8900
rect 44361 8851 44419 8857
rect 44836 8860 45928 8888
rect 31205 8823 31263 8829
rect 31205 8820 31217 8823
rect 28000 8792 31217 8820
rect 21453 8783 21511 8789
rect 31205 8789 31217 8792
rect 31251 8820 31263 8823
rect 31386 8820 31392 8832
rect 31251 8792 31392 8820
rect 31251 8789 31263 8792
rect 31205 8783 31263 8789
rect 31386 8780 31392 8792
rect 31444 8780 31450 8832
rect 32306 8780 32312 8832
rect 32364 8820 32370 8832
rect 34149 8823 34207 8829
rect 34149 8820 34161 8823
rect 32364 8792 34161 8820
rect 32364 8780 32370 8792
rect 34149 8789 34161 8792
rect 34195 8789 34207 8823
rect 34149 8783 34207 8789
rect 34238 8780 34244 8832
rect 34296 8820 34302 8832
rect 34977 8823 35035 8829
rect 34977 8820 34989 8823
rect 34296 8792 34989 8820
rect 34296 8780 34302 8792
rect 34977 8789 34989 8792
rect 35023 8789 35035 8823
rect 34977 8783 35035 8789
rect 35066 8780 35072 8832
rect 35124 8820 35130 8832
rect 36265 8823 36323 8829
rect 36265 8820 36277 8823
rect 35124 8792 36277 8820
rect 35124 8780 35130 8792
rect 36265 8789 36277 8792
rect 36311 8789 36323 8823
rect 36265 8783 36323 8789
rect 36633 8823 36691 8829
rect 36633 8789 36645 8823
rect 36679 8820 36691 8823
rect 36906 8820 36912 8832
rect 36679 8792 36912 8820
rect 36679 8789 36691 8792
rect 36633 8783 36691 8789
rect 36906 8780 36912 8792
rect 36964 8780 36970 8832
rect 37734 8780 37740 8832
rect 37792 8820 37798 8832
rect 38565 8823 38623 8829
rect 38565 8820 38577 8823
rect 37792 8792 38577 8820
rect 37792 8780 37798 8792
rect 38565 8789 38577 8792
rect 38611 8789 38623 8823
rect 38565 8783 38623 8789
rect 39114 8780 39120 8832
rect 39172 8820 39178 8832
rect 39853 8823 39911 8829
rect 39853 8820 39865 8823
rect 39172 8792 39865 8820
rect 39172 8780 39178 8792
rect 39853 8789 39865 8792
rect 39899 8789 39911 8823
rect 39853 8783 39911 8789
rect 42886 8780 42892 8832
rect 42944 8820 42950 8832
rect 44269 8823 44327 8829
rect 44269 8820 44281 8823
rect 42944 8792 44281 8820
rect 42944 8780 42950 8792
rect 44269 8789 44281 8792
rect 44315 8820 44327 8823
rect 44836 8820 44864 8860
rect 45922 8848 45928 8860
rect 45980 8848 45986 8900
rect 50172 8888 50200 8919
rect 50985 8891 51043 8897
rect 50985 8888 50997 8891
rect 46032 8860 50997 8888
rect 45186 8820 45192 8832
rect 44315 8792 44864 8820
rect 45147 8792 45192 8820
rect 44315 8789 44327 8792
rect 44269 8783 44327 8789
rect 45186 8780 45192 8792
rect 45244 8780 45250 8832
rect 45370 8780 45376 8832
rect 45428 8820 45434 8832
rect 46032 8820 46060 8860
rect 50985 8857 50997 8860
rect 51031 8888 51043 8891
rect 51031 8860 55812 8888
rect 51031 8857 51043 8860
rect 50985 8851 51043 8857
rect 45428 8792 46060 8820
rect 46293 8823 46351 8829
rect 45428 8780 45434 8792
rect 46293 8789 46305 8823
rect 46339 8820 46351 8823
rect 46382 8820 46388 8832
rect 46339 8792 46388 8820
rect 46339 8789 46351 8792
rect 46293 8783 46351 8789
rect 46382 8780 46388 8792
rect 46440 8820 46446 8832
rect 47670 8820 47676 8832
rect 46440 8792 47676 8820
rect 46440 8780 46446 8792
rect 47670 8780 47676 8792
rect 47728 8780 47734 8832
rect 55582 8820 55588 8832
rect 55543 8792 55588 8820
rect 55582 8780 55588 8792
rect 55640 8780 55646 8832
rect 55784 8820 55812 8860
rect 56594 8848 56600 8900
rect 56652 8848 56658 8900
rect 57790 8820 57796 8832
rect 55784 8792 57796 8820
rect 57790 8780 57796 8792
rect 57848 8780 57854 8832
rect 1104 8730 58880 8752
rect 1104 8678 15398 8730
rect 15450 8678 15462 8730
rect 15514 8678 15526 8730
rect 15578 8678 15590 8730
rect 15642 8678 15654 8730
rect 15706 8678 29846 8730
rect 29898 8678 29910 8730
rect 29962 8678 29974 8730
rect 30026 8678 30038 8730
rect 30090 8678 30102 8730
rect 30154 8678 44294 8730
rect 44346 8678 44358 8730
rect 44410 8678 44422 8730
rect 44474 8678 44486 8730
rect 44538 8678 44550 8730
rect 44602 8678 58880 8730
rect 1104 8656 58880 8678
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 17184 8588 18705 8616
rect 17184 8576 17190 8588
rect 18693 8585 18705 8588
rect 18739 8616 18751 8619
rect 19978 8616 19984 8628
rect 18739 8588 19984 8616
rect 18739 8585 18751 8588
rect 18693 8579 18751 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 26418 8576 26424 8628
rect 26476 8616 26482 8628
rect 28718 8616 28724 8628
rect 26476 8588 28724 8616
rect 26476 8576 26482 8588
rect 28718 8576 28724 8588
rect 28776 8576 28782 8628
rect 28813 8619 28871 8625
rect 28813 8585 28825 8619
rect 28859 8585 28871 8619
rect 29362 8616 29368 8628
rect 29323 8588 29368 8616
rect 28813 8579 28871 8585
rect 19889 8551 19947 8557
rect 19889 8517 19901 8551
rect 19935 8548 19947 8551
rect 20254 8548 20260 8560
rect 19935 8520 20260 8548
rect 19935 8517 19947 8520
rect 19889 8511 19947 8517
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 27341 8551 27399 8557
rect 27341 8548 27353 8551
rect 20364 8520 27353 8548
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 20364 8480 20392 8520
rect 27341 8517 27353 8520
rect 27387 8548 27399 8551
rect 27893 8551 27951 8557
rect 27893 8548 27905 8551
rect 27387 8520 27905 8548
rect 27387 8517 27399 8520
rect 27341 8511 27399 8517
rect 27893 8517 27905 8520
rect 27939 8548 27951 8551
rect 28166 8548 28172 8560
rect 27939 8520 28172 8548
rect 27939 8517 27951 8520
rect 27893 8511 27951 8517
rect 28166 8508 28172 8520
rect 28224 8548 28230 8560
rect 28828 8548 28856 8579
rect 29362 8576 29368 8588
rect 29420 8576 29426 8628
rect 29638 8576 29644 8628
rect 29696 8616 29702 8628
rect 30377 8619 30435 8625
rect 30377 8616 30389 8619
rect 29696 8588 30389 8616
rect 29696 8576 29702 8588
rect 30377 8585 30389 8588
rect 30423 8585 30435 8619
rect 31478 8616 31484 8628
rect 31439 8588 31484 8616
rect 30377 8579 30435 8585
rect 31478 8576 31484 8588
rect 31536 8576 31542 8628
rect 32674 8616 32680 8628
rect 32635 8588 32680 8616
rect 32674 8576 32680 8588
rect 32732 8576 32738 8628
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 33042 8616 33048 8628
rect 32824 8588 33048 8616
rect 32824 8576 32830 8588
rect 33042 8576 33048 8588
rect 33100 8616 33106 8628
rect 33459 8619 33517 8625
rect 33459 8616 33471 8619
rect 33100 8588 33471 8616
rect 33100 8576 33106 8588
rect 33459 8585 33471 8588
rect 33505 8585 33517 8619
rect 33459 8579 33517 8585
rect 34330 8576 34336 8628
rect 34388 8616 34394 8628
rect 35986 8616 35992 8628
rect 34388 8588 35992 8616
rect 34388 8576 34394 8588
rect 32122 8548 32128 8560
rect 28224 8520 28580 8548
rect 28828 8520 32128 8548
rect 28224 8508 28230 8520
rect 18840 8452 20392 8480
rect 20993 8483 21051 8489
rect 18840 8440 18846 8452
rect 20993 8449 21005 8483
rect 21039 8449 21051 8483
rect 28442 8480 28448 8492
rect 28403 8452 28448 8480
rect 20993 8443 21051 8449
rect 20349 8415 20407 8421
rect 20349 8381 20361 8415
rect 20395 8412 20407 8415
rect 21008 8412 21036 8443
rect 28442 8440 28448 8452
rect 28500 8440 28506 8492
rect 28552 8480 28580 8520
rect 29273 8483 29331 8489
rect 29273 8480 29285 8483
rect 28552 8452 29285 8480
rect 29273 8449 29285 8452
rect 29319 8449 29331 8483
rect 29273 8443 29331 8449
rect 29457 8483 29515 8489
rect 29457 8449 29469 8483
rect 29503 8480 29515 8483
rect 30282 8480 30288 8492
rect 29503 8452 30288 8480
rect 29503 8449 29515 8452
rect 29457 8443 29515 8449
rect 20395 8384 21036 8412
rect 28537 8415 28595 8421
rect 20395 8381 20407 8384
rect 20349 8375 20407 8381
rect 28537 8381 28549 8415
rect 28583 8381 28595 8415
rect 29288 8412 29316 8443
rect 30282 8440 30288 8452
rect 30340 8440 30346 8492
rect 30668 8489 30696 8520
rect 32122 8508 32128 8520
rect 32180 8508 32186 8560
rect 34624 8548 34652 8588
rect 35986 8576 35992 8588
rect 36044 8576 36050 8628
rect 36357 8619 36415 8625
rect 36357 8585 36369 8619
rect 36403 8616 36415 8619
rect 38470 8616 38476 8628
rect 36403 8588 38476 8616
rect 36403 8585 36415 8588
rect 36357 8579 36415 8585
rect 38470 8576 38476 8588
rect 38528 8576 38534 8628
rect 39942 8576 39948 8628
rect 40000 8616 40006 8628
rect 40954 8616 40960 8628
rect 40000 8588 40816 8616
rect 40915 8588 40960 8616
rect 40000 8576 40006 8588
rect 34546 8520 34652 8548
rect 35434 8508 35440 8560
rect 35492 8548 35498 8560
rect 39114 8548 39120 8560
rect 35492 8520 39120 8548
rect 35492 8508 35498 8520
rect 30561 8483 30619 8489
rect 30561 8449 30573 8483
rect 30607 8449 30619 8483
rect 30561 8443 30619 8449
rect 30653 8483 30711 8489
rect 30653 8449 30665 8483
rect 30699 8449 30711 8483
rect 30834 8480 30840 8492
rect 30795 8452 30840 8480
rect 30653 8443 30711 8449
rect 29288 8384 30420 8412
rect 28537 8375 28595 8381
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 20165 8347 20223 8353
rect 20165 8344 20177 8347
rect 20036 8316 20177 8344
rect 20036 8304 20042 8316
rect 20165 8313 20177 8316
rect 20211 8344 20223 8347
rect 20211 8316 20484 8344
rect 20211 8313 20223 8316
rect 20165 8307 20223 8313
rect 20456 8276 20484 8316
rect 20530 8304 20536 8356
rect 20588 8344 20594 8356
rect 20809 8347 20867 8353
rect 20809 8344 20821 8347
rect 20588 8316 20821 8344
rect 20588 8304 20594 8316
rect 20809 8313 20821 8316
rect 20855 8313 20867 8347
rect 28552 8344 28580 8375
rect 29638 8344 29644 8356
rect 28552 8316 29644 8344
rect 20809 8307 20867 8313
rect 29638 8304 29644 8316
rect 29696 8304 29702 8356
rect 21174 8276 21180 8288
rect 20456 8248 21180 8276
rect 21174 8236 21180 8248
rect 21232 8236 21238 8288
rect 27706 8236 27712 8288
rect 27764 8276 27770 8288
rect 28445 8279 28503 8285
rect 28445 8276 28457 8279
rect 27764 8248 28457 8276
rect 27764 8236 27770 8248
rect 28445 8245 28457 8248
rect 28491 8276 28503 8279
rect 28810 8276 28816 8288
rect 28491 8248 28816 8276
rect 28491 8245 28503 8248
rect 28445 8239 28503 8245
rect 28810 8236 28816 8248
rect 28868 8236 28874 8288
rect 30392 8276 30420 8384
rect 30466 8304 30472 8356
rect 30524 8344 30530 8356
rect 30576 8344 30604 8443
rect 30834 8440 30840 8452
rect 30892 8440 30898 8492
rect 30926 8440 30932 8492
rect 30984 8480 30990 8492
rect 32306 8480 32312 8492
rect 30984 8452 31029 8480
rect 31128 8452 32312 8480
rect 30984 8440 30990 8452
rect 30742 8372 30748 8424
rect 30800 8412 30806 8424
rect 31128 8412 31156 8452
rect 32306 8440 32312 8452
rect 32364 8440 32370 8492
rect 36280 8489 36308 8520
rect 39114 8508 39120 8520
rect 39172 8508 39178 8560
rect 39298 8508 39304 8560
rect 39356 8548 39362 8560
rect 39356 8520 40724 8548
rect 39356 8508 39362 8520
rect 35253 8483 35311 8489
rect 35253 8480 35265 8483
rect 34808 8452 35265 8480
rect 32030 8412 32036 8424
rect 30800 8384 31156 8412
rect 31220 8384 32036 8412
rect 30800 8372 30806 8384
rect 31220 8344 31248 8384
rect 32030 8372 32036 8384
rect 32088 8372 32094 8424
rect 32214 8412 32220 8424
rect 32175 8384 32220 8412
rect 32214 8372 32220 8384
rect 32272 8372 32278 8424
rect 32398 8372 32404 8424
rect 32456 8412 32462 8424
rect 34808 8412 34836 8452
rect 35253 8449 35265 8452
rect 35299 8449 35311 8483
rect 35253 8443 35311 8449
rect 36265 8483 36323 8489
rect 36265 8449 36277 8483
rect 36311 8449 36323 8483
rect 36265 8443 36323 8449
rect 36541 8483 36599 8489
rect 36541 8449 36553 8483
rect 36587 8449 36599 8483
rect 36541 8443 36599 8449
rect 32456 8384 34836 8412
rect 32456 8372 32462 8384
rect 34882 8372 34888 8424
rect 34940 8412 34946 8424
rect 34940 8384 34985 8412
rect 34940 8372 34946 8384
rect 31754 8344 31760 8356
rect 30524 8316 31248 8344
rect 31312 8316 31760 8344
rect 30524 8304 30530 8316
rect 31312 8276 31340 8316
rect 31754 8304 31760 8316
rect 31812 8304 31818 8356
rect 35805 8347 35863 8353
rect 35805 8313 35817 8347
rect 35851 8344 35863 8347
rect 36556 8344 36584 8443
rect 36906 8440 36912 8492
rect 36964 8480 36970 8492
rect 38562 8489 38568 8492
rect 37461 8483 37519 8489
rect 37461 8480 37473 8483
rect 36964 8452 37473 8480
rect 36964 8440 36970 8452
rect 37461 8449 37473 8452
rect 37507 8449 37519 8483
rect 38551 8483 38568 8489
rect 37461 8443 37519 8449
rect 37568 8452 38516 8480
rect 36725 8415 36783 8421
rect 36725 8381 36737 8415
rect 36771 8412 36783 8415
rect 37369 8415 37427 8421
rect 37369 8412 37381 8415
rect 36771 8384 37381 8412
rect 36771 8381 36783 8384
rect 36725 8375 36783 8381
rect 37369 8381 37381 8384
rect 37415 8381 37427 8415
rect 37369 8375 37427 8381
rect 37568 8344 37596 8452
rect 38378 8412 38384 8424
rect 38339 8384 38384 8412
rect 38378 8372 38384 8384
rect 38436 8372 38442 8424
rect 38488 8412 38516 8452
rect 38551 8449 38563 8483
rect 38551 8443 38568 8449
rect 38562 8440 38568 8443
rect 38620 8440 38626 8492
rect 39850 8480 39856 8492
rect 39811 8452 39856 8480
rect 39850 8440 39856 8452
rect 39908 8440 39914 8492
rect 40696 8489 40724 8520
rect 40788 8489 40816 8588
rect 40954 8576 40960 8588
rect 41012 8576 41018 8628
rect 42429 8619 42487 8625
rect 42429 8616 42441 8619
rect 41064 8588 42441 8616
rect 41064 8548 41092 8588
rect 42429 8585 42441 8588
rect 42475 8616 42487 8619
rect 42886 8616 42892 8628
rect 42475 8588 42892 8616
rect 42475 8585 42487 8588
rect 42429 8579 42487 8585
rect 42886 8576 42892 8588
rect 42944 8576 42950 8628
rect 44726 8616 44732 8628
rect 43180 8588 44732 8616
rect 43180 8557 43208 8588
rect 44726 8576 44732 8588
rect 44784 8576 44790 8628
rect 45094 8576 45100 8628
rect 45152 8616 45158 8628
rect 45281 8619 45339 8625
rect 45281 8616 45293 8619
rect 45152 8588 45293 8616
rect 45152 8576 45158 8588
rect 45281 8585 45293 8588
rect 45327 8585 45339 8619
rect 45281 8579 45339 8585
rect 45465 8619 45523 8625
rect 45465 8585 45477 8619
rect 45511 8616 45523 8619
rect 45554 8616 45560 8628
rect 45511 8588 45560 8616
rect 45511 8585 45523 8588
rect 45465 8579 45523 8585
rect 45554 8576 45560 8588
rect 45612 8576 45618 8628
rect 46198 8616 46204 8628
rect 46159 8588 46204 8616
rect 46198 8576 46204 8588
rect 46256 8576 46262 8628
rect 55398 8616 55404 8628
rect 55359 8588 55404 8616
rect 55398 8576 55404 8588
rect 55456 8576 55462 8628
rect 40880 8520 41092 8548
rect 43165 8551 43223 8557
rect 40681 8483 40739 8489
rect 40681 8449 40693 8483
rect 40727 8449 40739 8483
rect 40681 8443 40739 8449
rect 40773 8483 40831 8489
rect 40773 8449 40785 8483
rect 40819 8449 40831 8483
rect 40773 8443 40831 8449
rect 39666 8412 39672 8424
rect 38488 8384 39672 8412
rect 39666 8372 39672 8384
rect 39724 8372 39730 8424
rect 39942 8372 39948 8424
rect 40000 8412 40006 8424
rect 40880 8412 40908 8520
rect 43165 8517 43177 8551
rect 43211 8517 43223 8551
rect 45649 8551 45707 8557
rect 45649 8548 45661 8551
rect 43165 8511 43223 8517
rect 44376 8520 45661 8548
rect 44376 8492 44404 8520
rect 45649 8517 45661 8520
rect 45695 8517 45707 8551
rect 45649 8511 45707 8517
rect 41598 8480 41604 8492
rect 41559 8452 41604 8480
rect 41598 8440 41604 8452
rect 41656 8440 41662 8492
rect 44358 8480 44364 8492
rect 44319 8452 44364 8480
rect 44358 8440 44364 8452
rect 44416 8440 44422 8492
rect 44634 8480 44640 8492
rect 44595 8452 44640 8480
rect 44634 8440 44640 8452
rect 44692 8480 44698 8492
rect 45094 8480 45100 8492
rect 44692 8452 45100 8480
rect 44692 8440 44698 8452
rect 45094 8440 45100 8452
rect 45152 8440 45158 8492
rect 45370 8480 45376 8492
rect 45331 8452 45376 8480
rect 45370 8440 45376 8452
rect 45428 8440 45434 8492
rect 46382 8480 46388 8492
rect 46343 8452 46388 8480
rect 46382 8440 46388 8452
rect 46440 8440 46446 8492
rect 46566 8480 46572 8492
rect 46527 8452 46572 8480
rect 46566 8440 46572 8452
rect 46624 8440 46630 8492
rect 46661 8483 46719 8489
rect 46661 8449 46673 8483
rect 46707 8480 46719 8483
rect 47302 8480 47308 8492
rect 46707 8452 47308 8480
rect 46707 8449 46719 8452
rect 46661 8443 46719 8449
rect 47302 8440 47308 8452
rect 47360 8440 47366 8492
rect 40000 8384 40908 8412
rect 40000 8372 40006 8384
rect 40954 8372 40960 8424
rect 41012 8412 41018 8424
rect 41012 8384 41057 8412
rect 41012 8372 41018 8384
rect 42610 8372 42616 8424
rect 42668 8412 42674 8424
rect 44545 8415 44603 8421
rect 42668 8384 44312 8412
rect 42668 8372 42674 8384
rect 35851 8316 37596 8344
rect 37829 8347 37887 8353
rect 35851 8313 35863 8316
rect 35805 8307 35863 8313
rect 37829 8313 37841 8347
rect 37875 8344 37887 8347
rect 38470 8344 38476 8356
rect 37875 8316 38476 8344
rect 37875 8313 37887 8316
rect 37829 8307 37887 8313
rect 30392 8248 31340 8276
rect 31570 8236 31576 8288
rect 31628 8276 31634 8288
rect 34146 8276 34152 8288
rect 31628 8248 34152 8276
rect 31628 8236 31634 8248
rect 34146 8236 34152 8248
rect 34204 8236 34210 8288
rect 34514 8236 34520 8288
rect 34572 8276 34578 8288
rect 35820 8276 35848 8307
rect 38470 8304 38476 8316
rect 38528 8304 38534 8356
rect 38841 8347 38899 8353
rect 38841 8313 38853 8347
rect 38887 8344 38899 8347
rect 39758 8344 39764 8356
rect 38887 8316 39764 8344
rect 38887 8313 38899 8316
rect 38841 8307 38899 8313
rect 39758 8304 39764 8316
rect 39816 8304 39822 8356
rect 41414 8304 41420 8356
rect 41472 8344 41478 8356
rect 44177 8347 44235 8353
rect 44177 8344 44189 8347
rect 41472 8316 41517 8344
rect 42352 8316 44189 8344
rect 41472 8304 41478 8316
rect 34572 8248 35848 8276
rect 34572 8236 34578 8248
rect 37458 8236 37464 8288
rect 37516 8276 37522 8288
rect 39942 8276 39948 8288
rect 37516 8248 39948 8276
rect 37516 8236 37522 8248
rect 39942 8236 39948 8248
rect 40000 8236 40006 8288
rect 40221 8279 40279 8285
rect 40221 8245 40233 8279
rect 40267 8276 40279 8279
rect 40402 8276 40408 8288
rect 40267 8248 40408 8276
rect 40267 8245 40279 8248
rect 40221 8239 40279 8245
rect 40402 8236 40408 8248
rect 40460 8236 40466 8288
rect 40494 8236 40500 8288
rect 40552 8276 40558 8288
rect 41322 8276 41328 8288
rect 40552 8248 41328 8276
rect 40552 8236 40558 8248
rect 41322 8236 41328 8248
rect 41380 8276 41386 8288
rect 42352 8276 42380 8316
rect 44177 8313 44189 8316
rect 44223 8313 44235 8347
rect 44284 8344 44312 8384
rect 44545 8381 44557 8415
rect 44591 8412 44603 8415
rect 45388 8412 45416 8440
rect 44591 8384 45416 8412
rect 44591 8381 44603 8384
rect 44545 8375 44603 8381
rect 45097 8347 45155 8353
rect 45097 8344 45109 8347
rect 44284 8316 45109 8344
rect 44177 8307 44235 8313
rect 45097 8313 45109 8316
rect 45143 8313 45155 8347
rect 45097 8307 45155 8313
rect 43070 8276 43076 8288
rect 41380 8248 42380 8276
rect 43031 8248 43076 8276
rect 41380 8236 41386 8248
rect 43070 8236 43076 8248
rect 43128 8236 43134 8288
rect 44266 8236 44272 8288
rect 44324 8276 44330 8288
rect 44361 8279 44419 8285
rect 44361 8276 44373 8279
rect 44324 8248 44373 8276
rect 44324 8236 44330 8248
rect 44361 8245 44373 8248
rect 44407 8245 44419 8279
rect 44361 8239 44419 8245
rect 1104 8186 58880 8208
rect 1104 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 8302 8186
rect 8354 8134 8366 8186
rect 8418 8134 8430 8186
rect 8482 8134 22622 8186
rect 22674 8134 22686 8186
rect 22738 8134 22750 8186
rect 22802 8134 22814 8186
rect 22866 8134 22878 8186
rect 22930 8134 37070 8186
rect 37122 8134 37134 8186
rect 37186 8134 37198 8186
rect 37250 8134 37262 8186
rect 37314 8134 37326 8186
rect 37378 8134 51518 8186
rect 51570 8134 51582 8186
rect 51634 8134 51646 8186
rect 51698 8134 51710 8186
rect 51762 8134 51774 8186
rect 51826 8134 58880 8186
rect 1104 8112 58880 8134
rect 21174 8072 21180 8084
rect 21135 8044 21180 8072
rect 21174 8032 21180 8044
rect 21232 8032 21238 8084
rect 26418 8032 26424 8084
rect 26476 8072 26482 8084
rect 26881 8075 26939 8081
rect 26881 8072 26893 8075
rect 26476 8044 26893 8072
rect 26476 8032 26482 8044
rect 26881 8041 26893 8044
rect 26927 8041 26939 8075
rect 26881 8035 26939 8041
rect 28077 8075 28135 8081
rect 28077 8041 28089 8075
rect 28123 8072 28135 8075
rect 28166 8072 28172 8084
rect 28123 8044 28172 8072
rect 28123 8041 28135 8044
rect 28077 8035 28135 8041
rect 28166 8032 28172 8044
rect 28224 8032 28230 8084
rect 30834 8072 30840 8084
rect 30795 8044 30840 8072
rect 30834 8032 30840 8044
rect 30892 8032 30898 8084
rect 32214 8032 32220 8084
rect 32272 8072 32278 8084
rect 32769 8075 32827 8081
rect 32769 8072 32781 8075
rect 32272 8044 32781 8072
rect 32272 8032 32278 8044
rect 32769 8041 32781 8044
rect 32815 8041 32827 8075
rect 32769 8035 32827 8041
rect 33042 8032 33048 8084
rect 33100 8072 33106 8084
rect 33100 8044 36032 8072
rect 33100 8032 33106 8044
rect 29825 8007 29883 8013
rect 29825 7973 29837 8007
rect 29871 8004 29883 8007
rect 30926 8004 30932 8016
rect 29871 7976 30932 8004
rect 29871 7973 29883 7976
rect 29825 7967 29883 7973
rect 30926 7964 30932 7976
rect 30984 7964 30990 8016
rect 31662 8004 31668 8016
rect 31623 7976 31668 8004
rect 31662 7964 31668 7976
rect 31720 7964 31726 8016
rect 31754 7964 31760 8016
rect 31812 8004 31818 8016
rect 36004 8004 36032 8044
rect 36906 8032 36912 8084
rect 36964 8072 36970 8084
rect 37001 8075 37059 8081
rect 37001 8072 37013 8075
rect 36964 8044 37013 8072
rect 36964 8032 36970 8044
rect 37001 8041 37013 8044
rect 37047 8041 37059 8075
rect 40218 8072 40224 8084
rect 37001 8035 37059 8041
rect 38764 8044 40224 8072
rect 37458 8004 37464 8016
rect 31812 7976 34836 8004
rect 36004 7976 37464 8004
rect 31812 7964 31818 7976
rect 27798 7896 27804 7948
rect 27856 7936 27862 7948
rect 27893 7939 27951 7945
rect 27893 7936 27905 7939
rect 27856 7908 27905 7936
rect 27856 7896 27862 7908
rect 27893 7905 27905 7908
rect 27939 7936 27951 7939
rect 28626 7936 28632 7948
rect 27939 7908 28632 7936
rect 27939 7905 27951 7908
rect 27893 7899 27951 7905
rect 28626 7896 28632 7908
rect 28684 7896 28690 7948
rect 28997 7939 29055 7945
rect 28997 7905 29009 7939
rect 29043 7936 29055 7939
rect 29454 7936 29460 7948
rect 29043 7908 29460 7936
rect 29043 7905 29055 7908
rect 28997 7899 29055 7905
rect 29454 7896 29460 7908
rect 29512 7896 29518 7948
rect 30558 7936 30564 7948
rect 30519 7908 30564 7936
rect 30558 7896 30564 7908
rect 30616 7896 30622 7948
rect 32214 7936 32220 7948
rect 31726 7908 32220 7936
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 20438 7868 20444 7880
rect 20395 7840 20444 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 28074 7868 28080 7880
rect 20588 7840 20633 7868
rect 28035 7840 28080 7868
rect 20588 7828 20594 7840
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 28718 7868 28724 7880
rect 28679 7840 28724 7868
rect 28718 7828 28724 7840
rect 28776 7828 28782 7880
rect 28813 7871 28871 7877
rect 28813 7837 28825 7871
rect 28859 7868 28871 7871
rect 29730 7868 29736 7880
rect 28859 7840 29736 7868
rect 28859 7837 28871 7840
rect 28813 7831 28871 7837
rect 29730 7828 29736 7840
rect 29788 7828 29794 7880
rect 30469 7871 30527 7877
rect 30469 7837 30481 7871
rect 30515 7868 30527 7871
rect 31726 7868 31754 7908
rect 32214 7896 32220 7908
rect 32272 7936 32278 7948
rect 33042 7936 33048 7948
rect 32272 7908 33048 7936
rect 32272 7896 32278 7908
rect 33042 7896 33048 7908
rect 33100 7896 33106 7948
rect 34238 7936 34244 7948
rect 33704 7908 34244 7936
rect 33704 7880 33732 7908
rect 34238 7896 34244 7908
rect 34296 7896 34302 7948
rect 34698 7936 34704 7948
rect 34659 7908 34704 7936
rect 34698 7896 34704 7908
rect 34756 7896 34762 7948
rect 34808 7936 34836 7976
rect 37458 7964 37464 7976
rect 37516 7964 37522 8016
rect 36449 7939 36507 7945
rect 36449 7936 36461 7939
rect 34808 7908 36461 7936
rect 36449 7905 36461 7908
rect 36495 7905 36507 7939
rect 38470 7936 38476 7948
rect 38431 7908 38476 7936
rect 36449 7899 36507 7905
rect 38470 7896 38476 7908
rect 38528 7896 38534 7948
rect 38764 7945 38792 8044
rect 40218 8032 40224 8044
rect 40276 8032 40282 8084
rect 41877 8075 41935 8081
rect 41877 8041 41889 8075
rect 41923 8072 41935 8075
rect 44358 8072 44364 8084
rect 41923 8044 44364 8072
rect 41923 8041 41935 8044
rect 41877 8035 41935 8041
rect 44358 8032 44364 8044
rect 44416 8032 44422 8084
rect 47302 8072 47308 8084
rect 47263 8044 47308 8072
rect 47302 8032 47308 8044
rect 47360 8032 47366 8084
rect 39301 8007 39359 8013
rect 39301 7973 39313 8007
rect 39347 8004 39359 8007
rect 39850 8004 39856 8016
rect 39347 7976 39856 8004
rect 39347 7973 39359 7976
rect 39301 7967 39359 7973
rect 39850 7964 39856 7976
rect 39908 7964 39914 8016
rect 45005 8007 45063 8013
rect 45005 7973 45017 8007
rect 45051 7973 45063 8007
rect 45005 7967 45063 7973
rect 38749 7939 38807 7945
rect 38749 7905 38761 7939
rect 38795 7905 38807 7939
rect 38749 7899 38807 7905
rect 40034 7896 40040 7948
rect 40092 7936 40098 7948
rect 40129 7939 40187 7945
rect 40129 7936 40141 7939
rect 40092 7908 40141 7936
rect 40092 7896 40098 7908
rect 40129 7905 40141 7908
rect 40175 7936 40187 7939
rect 42334 7936 42340 7948
rect 40175 7908 42340 7936
rect 40175 7905 40187 7908
rect 40129 7899 40187 7905
rect 42334 7896 42340 7908
rect 42392 7896 42398 7948
rect 42613 7939 42671 7945
rect 42613 7905 42625 7939
rect 42659 7936 42671 7939
rect 45020 7936 45048 7967
rect 57790 7964 57796 8016
rect 57848 8004 57854 8016
rect 57885 8007 57943 8013
rect 57885 8004 57897 8007
rect 57848 7976 57897 8004
rect 57848 7964 57854 7976
rect 57885 7973 57897 7976
rect 57931 7973 57943 8007
rect 57885 7967 57943 7973
rect 42659 7908 45048 7936
rect 45465 7939 45523 7945
rect 42659 7905 42671 7908
rect 42613 7899 42671 7905
rect 45465 7905 45477 7939
rect 45511 7936 45523 7939
rect 46017 7939 46075 7945
rect 46017 7936 46029 7939
rect 45511 7908 46029 7936
rect 45511 7905 45523 7908
rect 45465 7899 45523 7905
rect 46017 7905 46029 7908
rect 46063 7905 46075 7939
rect 46382 7936 46388 7948
rect 46017 7899 46075 7905
rect 46216 7908 46388 7936
rect 30515 7840 31754 7868
rect 30515 7837 30527 7840
rect 30469 7831 30527 7837
rect 32030 7828 32036 7880
rect 32088 7868 32094 7880
rect 32309 7871 32367 7877
rect 32309 7868 32321 7871
rect 32088 7840 32321 7868
rect 32088 7828 32094 7840
rect 32309 7837 32321 7840
rect 32355 7837 32367 7871
rect 32309 7831 32367 7837
rect 32490 7828 32496 7880
rect 32548 7868 32554 7880
rect 32585 7871 32643 7877
rect 32585 7868 32597 7871
rect 32548 7840 32597 7868
rect 32548 7828 32554 7840
rect 32585 7837 32597 7840
rect 32631 7837 32643 7871
rect 33686 7868 33692 7880
rect 33599 7840 33692 7868
rect 32585 7831 32643 7837
rect 33686 7828 33692 7840
rect 33744 7828 33750 7880
rect 33965 7871 34023 7877
rect 33965 7837 33977 7871
rect 34011 7868 34023 7871
rect 34514 7868 34520 7880
rect 34011 7840 34520 7868
rect 34011 7837 34023 7840
rect 33965 7831 34023 7837
rect 34514 7828 34520 7840
rect 34572 7828 34578 7880
rect 45370 7868 45376 7880
rect 45283 7840 45376 7868
rect 45370 7828 45376 7840
rect 45428 7828 45434 7880
rect 46216 7877 46244 7908
rect 46382 7896 46388 7908
rect 46440 7896 46446 7948
rect 46201 7871 46259 7877
rect 46201 7837 46213 7871
rect 46247 7837 46259 7871
rect 46201 7831 46259 7837
rect 46290 7828 46296 7880
rect 46348 7868 46354 7880
rect 46477 7871 46535 7877
rect 46477 7868 46489 7871
rect 46348 7840 46489 7868
rect 46348 7828 46354 7840
rect 46477 7837 46489 7840
rect 46523 7868 46535 7871
rect 46937 7871 46995 7877
rect 46937 7868 46949 7871
rect 46523 7840 46949 7868
rect 46523 7837 46535 7840
rect 46477 7831 46535 7837
rect 46937 7837 46949 7840
rect 46983 7837 46995 7871
rect 46937 7831 46995 7837
rect 27798 7800 27804 7812
rect 27759 7772 27804 7800
rect 27798 7760 27804 7772
rect 27856 7760 27862 7812
rect 28997 7803 29055 7809
rect 28997 7769 29009 7803
rect 29043 7800 29055 7803
rect 31294 7800 31300 7812
rect 29043 7772 31300 7800
rect 29043 7769 29055 7772
rect 28997 7763 29055 7769
rect 31294 7760 31300 7772
rect 31352 7760 31358 7812
rect 31389 7803 31447 7809
rect 31389 7769 31401 7803
rect 31435 7800 31447 7803
rect 31570 7800 31576 7812
rect 31435 7772 31576 7800
rect 31435 7769 31447 7772
rect 31389 7763 31447 7769
rect 20717 7735 20775 7741
rect 20717 7701 20729 7735
rect 20763 7732 20775 7735
rect 20898 7732 20904 7744
rect 20763 7704 20904 7732
rect 20763 7701 20775 7704
rect 20717 7695 20775 7701
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 28261 7735 28319 7741
rect 28261 7701 28273 7735
rect 28307 7732 28319 7735
rect 28442 7732 28448 7744
rect 28307 7704 28448 7732
rect 28307 7701 28319 7704
rect 28261 7695 28319 7701
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 29086 7692 29092 7744
rect 29144 7732 29150 7744
rect 31404 7732 31432 7763
rect 31570 7760 31576 7772
rect 31628 7760 31634 7812
rect 32122 7760 32128 7812
rect 32180 7800 32186 7812
rect 32401 7803 32459 7809
rect 32401 7800 32413 7803
rect 32180 7772 32413 7800
rect 32180 7760 32186 7772
rect 32401 7769 32413 7772
rect 32447 7769 32459 7803
rect 32401 7763 32459 7769
rect 32674 7760 32680 7812
rect 32732 7800 32738 7812
rect 34977 7803 35035 7809
rect 34977 7800 34989 7803
rect 32732 7772 34989 7800
rect 32732 7760 32738 7772
rect 34977 7769 34989 7772
rect 35023 7769 35035 7803
rect 34977 7763 35035 7769
rect 35986 7760 35992 7812
rect 36044 7760 36050 7812
rect 38010 7760 38016 7812
rect 38068 7800 38074 7812
rect 38470 7800 38476 7812
rect 38068 7772 38476 7800
rect 38068 7760 38074 7772
rect 38470 7760 38476 7772
rect 38528 7760 38534 7812
rect 40402 7800 40408 7812
rect 40363 7772 40408 7800
rect 40402 7760 40408 7772
rect 40460 7760 40466 7812
rect 41690 7800 41696 7812
rect 41630 7772 41696 7800
rect 41690 7760 41696 7772
rect 41748 7760 41754 7812
rect 43162 7760 43168 7812
rect 43220 7760 43226 7812
rect 45388 7800 45416 7828
rect 47118 7800 47124 7812
rect 44100 7772 47124 7800
rect 31846 7732 31852 7744
rect 29144 7704 31432 7732
rect 31807 7704 31852 7732
rect 29144 7692 29150 7704
rect 31846 7692 31852 7704
rect 31904 7692 31910 7744
rect 33778 7732 33784 7744
rect 33739 7704 33784 7732
rect 33778 7692 33784 7704
rect 33836 7692 33842 7744
rect 34149 7735 34207 7741
rect 34149 7701 34161 7735
rect 34195 7732 34207 7735
rect 34330 7732 34336 7744
rect 34195 7704 34336 7732
rect 34195 7701 34207 7704
rect 34149 7695 34207 7701
rect 34330 7692 34336 7704
rect 34388 7692 34394 7744
rect 44100 7741 44128 7772
rect 47118 7760 47124 7772
rect 47176 7760 47182 7812
rect 57425 7803 57483 7809
rect 57425 7769 57437 7803
rect 57471 7800 57483 7803
rect 58066 7800 58072 7812
rect 57471 7772 58072 7800
rect 57471 7769 57483 7772
rect 57425 7763 57483 7769
rect 58066 7760 58072 7772
rect 58124 7760 58130 7812
rect 44085 7735 44143 7741
rect 44085 7701 44097 7735
rect 44131 7701 44143 7735
rect 46382 7732 46388 7744
rect 46343 7704 46388 7732
rect 44085 7695 44143 7701
rect 46382 7692 46388 7704
rect 46440 7692 46446 7744
rect 1104 7642 58880 7664
rect 1104 7590 15398 7642
rect 15450 7590 15462 7642
rect 15514 7590 15526 7642
rect 15578 7590 15590 7642
rect 15642 7590 15654 7642
rect 15706 7590 29846 7642
rect 29898 7590 29910 7642
rect 29962 7590 29974 7642
rect 30026 7590 30038 7642
rect 30090 7590 30102 7642
rect 30154 7590 44294 7642
rect 44346 7590 44358 7642
rect 44410 7590 44422 7642
rect 44474 7590 44486 7642
rect 44538 7590 44550 7642
rect 44602 7590 58880 7642
rect 1104 7568 58880 7590
rect 27341 7531 27399 7537
rect 27341 7497 27353 7531
rect 27387 7528 27399 7531
rect 27614 7528 27620 7540
rect 27387 7500 27620 7528
rect 27387 7497 27399 7500
rect 27341 7491 27399 7497
rect 27614 7488 27620 7500
rect 27672 7528 27678 7540
rect 28074 7528 28080 7540
rect 27672 7500 28080 7528
rect 27672 7488 27678 7500
rect 28074 7488 28080 7500
rect 28132 7488 28138 7540
rect 28718 7488 28724 7540
rect 28776 7528 28782 7540
rect 28997 7531 29055 7537
rect 28997 7528 29009 7531
rect 28776 7500 29009 7528
rect 28776 7488 28782 7500
rect 28997 7497 29009 7500
rect 29043 7497 29055 7531
rect 28997 7491 29055 7497
rect 29730 7488 29736 7540
rect 29788 7528 29794 7540
rect 29917 7531 29975 7537
rect 29917 7528 29929 7531
rect 29788 7500 29929 7528
rect 29788 7488 29794 7500
rect 29917 7497 29929 7500
rect 29963 7497 29975 7531
rect 32674 7528 32680 7540
rect 32635 7500 32680 7528
rect 29917 7491 29975 7497
rect 32674 7488 32680 7500
rect 32732 7488 32738 7540
rect 34422 7528 34428 7540
rect 33704 7500 34428 7528
rect 7558 7420 7564 7472
rect 7616 7460 7622 7472
rect 21634 7460 21640 7472
rect 7616 7432 21640 7460
rect 7616 7420 7622 7432
rect 21634 7420 21640 7432
rect 21692 7460 21698 7472
rect 29178 7469 29184 7472
rect 22005 7463 22063 7469
rect 22005 7460 22017 7463
rect 21692 7432 22017 7460
rect 21692 7420 21698 7432
rect 22005 7429 22017 7432
rect 22051 7429 22063 7463
rect 22005 7423 22063 7429
rect 29165 7463 29184 7469
rect 29165 7429 29177 7463
rect 29165 7423 29184 7429
rect 29178 7420 29184 7423
rect 29236 7420 29242 7472
rect 33704 7469 33732 7500
rect 34422 7488 34428 7500
rect 34480 7488 34486 7540
rect 37645 7531 37703 7537
rect 37645 7497 37657 7531
rect 37691 7528 37703 7531
rect 38378 7528 38384 7540
rect 37691 7500 38384 7528
rect 37691 7497 37703 7500
rect 37645 7491 37703 7497
rect 38378 7488 38384 7500
rect 38436 7488 38442 7540
rect 38470 7488 38476 7540
rect 38528 7528 38534 7540
rect 38528 7500 40264 7528
rect 38528 7488 38534 7500
rect 29365 7463 29423 7469
rect 29365 7429 29377 7463
rect 29411 7429 29423 7463
rect 33505 7463 33563 7469
rect 33505 7460 33517 7463
rect 29365 7423 29423 7429
rect 31128 7432 33517 7460
rect 20898 7392 20904 7404
rect 20859 7364 20904 7392
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 27525 7395 27583 7401
rect 27525 7361 27537 7395
rect 27571 7392 27583 7395
rect 28258 7392 28264 7404
rect 27571 7364 28264 7392
rect 27571 7361 27583 7364
rect 27525 7355 27583 7361
rect 28258 7352 28264 7364
rect 28316 7352 28322 7404
rect 28626 7352 28632 7404
rect 28684 7392 28690 7404
rect 29380 7392 29408 7423
rect 28684 7364 29408 7392
rect 28684 7352 28690 7364
rect 29638 7352 29644 7404
rect 29696 7392 29702 7404
rect 29825 7395 29883 7401
rect 29825 7392 29837 7395
rect 29696 7364 29837 7392
rect 29696 7352 29702 7364
rect 29825 7361 29837 7364
rect 29871 7361 29883 7395
rect 29825 7355 29883 7361
rect 30009 7395 30067 7401
rect 30009 7361 30021 7395
rect 30055 7392 30067 7395
rect 30742 7392 30748 7404
rect 30055 7364 30748 7392
rect 30055 7361 30067 7364
rect 30009 7355 30067 7361
rect 21913 7327 21971 7333
rect 21913 7293 21925 7327
rect 21959 7293 21971 7327
rect 21913 7287 21971 7293
rect 21085 7259 21143 7265
rect 21085 7225 21097 7259
rect 21131 7256 21143 7259
rect 21928 7256 21956 7287
rect 27706 7284 27712 7336
rect 27764 7324 27770 7336
rect 28077 7327 28135 7333
rect 28077 7324 28089 7327
rect 27764 7296 28089 7324
rect 27764 7284 27770 7296
rect 28077 7293 28089 7296
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 28169 7327 28227 7333
rect 28169 7293 28181 7327
rect 28215 7293 28227 7327
rect 28350 7324 28356 7336
rect 28311 7296 28356 7324
rect 28169 7287 28227 7293
rect 21131 7228 21956 7256
rect 22465 7259 22523 7265
rect 21131 7225 21143 7228
rect 21085 7219 21143 7225
rect 22465 7225 22477 7259
rect 22511 7225 22523 7259
rect 22465 7219 22523 7225
rect 22480 7188 22508 7219
rect 27982 7216 27988 7268
rect 28040 7256 28046 7268
rect 28184 7256 28212 7287
rect 28350 7284 28356 7296
rect 28408 7284 28414 7336
rect 28442 7284 28448 7336
rect 28500 7324 28506 7336
rect 30024 7324 30052 7355
rect 30742 7352 30748 7364
rect 30800 7352 30806 7404
rect 31128 7401 31156 7432
rect 33505 7429 33517 7432
rect 33551 7429 33563 7463
rect 33505 7423 33563 7429
rect 33689 7463 33747 7469
rect 33689 7429 33701 7463
rect 33735 7429 33747 7463
rect 39408 7460 39436 7500
rect 39758 7460 39764 7472
rect 39330 7432 39436 7460
rect 39719 7432 39764 7460
rect 33689 7423 33747 7429
rect 39758 7420 39764 7432
rect 39816 7420 39822 7472
rect 31113 7395 31171 7401
rect 31113 7392 31125 7395
rect 30852 7364 31125 7392
rect 28500 7296 30052 7324
rect 28500 7284 28506 7296
rect 30852 7256 30880 7364
rect 31113 7361 31125 7364
rect 31159 7361 31171 7395
rect 31113 7355 31171 7361
rect 31570 7352 31576 7404
rect 31628 7392 31634 7404
rect 32309 7395 32367 7401
rect 32309 7392 32321 7395
rect 31628 7364 32321 7392
rect 31628 7352 31634 7364
rect 32309 7361 32321 7364
rect 32355 7361 32367 7395
rect 32309 7355 32367 7361
rect 33042 7352 33048 7404
rect 33100 7392 33106 7404
rect 34238 7392 34244 7404
rect 33100 7364 34244 7392
rect 33100 7352 33106 7364
rect 34238 7352 34244 7364
rect 34296 7392 34302 7404
rect 34425 7395 34483 7401
rect 34425 7392 34437 7395
rect 34296 7364 34437 7392
rect 34296 7352 34302 7364
rect 34425 7361 34437 7364
rect 34471 7361 34483 7395
rect 34425 7355 34483 7361
rect 37553 7395 37611 7401
rect 37553 7361 37565 7395
rect 37599 7361 37611 7395
rect 37734 7392 37740 7404
rect 37695 7364 37740 7392
rect 37553 7355 37611 7361
rect 31202 7324 31208 7336
rect 31163 7296 31208 7324
rect 31202 7284 31208 7296
rect 31260 7284 31266 7336
rect 31294 7284 31300 7336
rect 31352 7324 31358 7336
rect 32217 7327 32275 7333
rect 32217 7324 32229 7327
rect 31352 7296 32229 7324
rect 31352 7284 31358 7296
rect 32217 7293 32229 7296
rect 32263 7293 32275 7327
rect 34330 7324 34336 7336
rect 34291 7296 34336 7324
rect 32217 7287 32275 7293
rect 34330 7284 34336 7296
rect 34388 7284 34394 7336
rect 28040 7228 30880 7256
rect 31481 7259 31539 7265
rect 28040 7216 28046 7228
rect 31481 7225 31493 7259
rect 31527 7256 31539 7259
rect 33594 7256 33600 7268
rect 31527 7228 33600 7256
rect 31527 7225 31539 7228
rect 31481 7219 31539 7225
rect 33594 7216 33600 7228
rect 33652 7216 33658 7268
rect 36722 7256 36728 7268
rect 36635 7228 36728 7256
rect 36722 7216 36728 7228
rect 36780 7256 36786 7268
rect 37568 7256 37596 7355
rect 37734 7352 37740 7364
rect 37792 7352 37798 7404
rect 40034 7352 40040 7404
rect 40092 7392 40098 7404
rect 40236 7392 40264 7500
rect 41138 7488 41144 7540
rect 41196 7528 41202 7540
rect 41325 7531 41383 7537
rect 41325 7528 41337 7531
rect 41196 7500 41337 7528
rect 41196 7488 41202 7500
rect 41325 7497 41337 7500
rect 41371 7497 41383 7531
rect 41325 7491 41383 7497
rect 44177 7531 44235 7537
rect 44177 7497 44189 7531
rect 44223 7528 44235 7531
rect 44634 7528 44640 7540
rect 44223 7500 44640 7528
rect 44223 7497 44235 7500
rect 44177 7491 44235 7497
rect 44634 7488 44640 7500
rect 44692 7488 44698 7540
rect 44726 7488 44732 7540
rect 44784 7528 44790 7540
rect 46109 7531 46167 7537
rect 44784 7500 44829 7528
rect 44784 7488 44790 7500
rect 46109 7497 46121 7531
rect 46155 7528 46167 7531
rect 46290 7528 46296 7540
rect 46155 7500 46296 7528
rect 46155 7497 46167 7500
rect 46109 7491 46167 7497
rect 46290 7488 46296 7500
rect 46348 7488 46354 7540
rect 46566 7528 46572 7540
rect 46527 7500 46572 7528
rect 46566 7488 46572 7500
rect 46624 7488 46630 7540
rect 40402 7420 40408 7472
rect 40460 7460 40466 7472
rect 40773 7463 40831 7469
rect 40773 7460 40785 7463
rect 40460 7432 40785 7460
rect 40460 7420 40466 7432
rect 40773 7429 40785 7432
rect 40819 7460 40831 7463
rect 41690 7460 41696 7472
rect 40819 7432 41696 7460
rect 40819 7429 40831 7432
rect 40773 7423 40831 7429
rect 41690 7420 41696 7432
rect 41748 7460 41754 7472
rect 43162 7460 43168 7472
rect 41748 7432 43168 7460
rect 41748 7420 41754 7432
rect 43162 7420 43168 7432
rect 43220 7420 43226 7472
rect 45554 7420 45560 7472
rect 45612 7460 45618 7472
rect 45741 7463 45799 7469
rect 45741 7460 45753 7463
rect 45612 7432 45753 7460
rect 45612 7420 45618 7432
rect 45741 7429 45753 7432
rect 45787 7460 45799 7463
rect 46661 7463 46719 7469
rect 46661 7460 46673 7463
rect 45787 7432 46673 7460
rect 45787 7429 45799 7432
rect 45741 7423 45799 7429
rect 46661 7429 46673 7432
rect 46707 7429 46719 7463
rect 46661 7423 46719 7429
rect 46845 7463 46903 7469
rect 46845 7429 46857 7463
rect 46891 7460 46903 7463
rect 47118 7460 47124 7472
rect 46891 7432 47124 7460
rect 46891 7429 46903 7432
rect 46845 7423 46903 7429
rect 47118 7420 47124 7432
rect 47176 7420 47182 7472
rect 40589 7395 40647 7401
rect 40589 7392 40601 7395
rect 40092 7364 40137 7392
rect 40236 7364 40601 7392
rect 40092 7352 40098 7364
rect 40589 7361 40601 7364
rect 40635 7361 40647 7395
rect 40589 7355 40647 7361
rect 41322 7352 41328 7404
rect 41380 7392 41386 7404
rect 41417 7395 41475 7401
rect 41417 7392 41429 7395
rect 41380 7364 41429 7392
rect 41380 7352 41386 7364
rect 41417 7361 41429 7364
rect 41463 7361 41475 7395
rect 41417 7355 41475 7361
rect 42334 7352 42340 7404
rect 42392 7392 42398 7404
rect 42429 7395 42487 7401
rect 42429 7392 42441 7395
rect 42392 7364 42441 7392
rect 42392 7352 42398 7364
rect 42429 7361 42441 7364
rect 42475 7361 42487 7395
rect 42429 7355 42487 7361
rect 44637 7395 44695 7401
rect 44637 7361 44649 7395
rect 44683 7392 44695 7395
rect 45094 7392 45100 7404
rect 44683 7364 45100 7392
rect 44683 7361 44695 7364
rect 44637 7355 44695 7361
rect 45094 7352 45100 7364
rect 45152 7392 45158 7404
rect 45462 7392 45468 7404
rect 45152 7364 45468 7392
rect 45152 7352 45158 7364
rect 45462 7352 45468 7364
rect 45520 7352 45526 7404
rect 45922 7392 45928 7404
rect 45883 7364 45928 7392
rect 45922 7352 45928 7364
rect 45980 7392 45986 7404
rect 46569 7395 46627 7401
rect 46569 7392 46581 7395
rect 45980 7364 46581 7392
rect 45980 7352 45986 7364
rect 46569 7361 46581 7364
rect 46615 7361 46627 7395
rect 46569 7355 46627 7361
rect 38289 7327 38347 7333
rect 38289 7293 38301 7327
rect 38335 7324 38347 7327
rect 38562 7324 38568 7336
rect 38335 7296 38568 7324
rect 38335 7293 38347 7296
rect 38289 7287 38347 7293
rect 38562 7284 38568 7296
rect 38620 7284 38626 7336
rect 39206 7324 39212 7336
rect 38672 7296 39212 7324
rect 38672 7256 38700 7296
rect 39206 7284 39212 7296
rect 39264 7284 39270 7336
rect 42705 7327 42763 7333
rect 42705 7293 42717 7327
rect 42751 7324 42763 7327
rect 45186 7324 45192 7336
rect 42751 7296 45192 7324
rect 42751 7293 42763 7296
rect 42705 7287 42763 7293
rect 45186 7284 45192 7296
rect 45244 7284 45250 7336
rect 36780 7228 38700 7256
rect 36780 7216 36786 7228
rect 28074 7188 28080 7200
rect 22480 7160 28080 7188
rect 28074 7148 28080 7160
rect 28132 7148 28138 7200
rect 28537 7191 28595 7197
rect 28537 7157 28549 7191
rect 28583 7188 28595 7191
rect 29086 7188 29092 7200
rect 28583 7160 29092 7188
rect 28583 7157 28595 7160
rect 28537 7151 28595 7157
rect 29086 7148 29092 7160
rect 29144 7148 29150 7200
rect 29181 7191 29239 7197
rect 29181 7157 29193 7191
rect 29227 7188 29239 7191
rect 29638 7188 29644 7200
rect 29227 7160 29644 7188
rect 29227 7157 29239 7160
rect 29181 7151 29239 7157
rect 29638 7148 29644 7160
rect 29696 7148 29702 7200
rect 34698 7188 34704 7200
rect 34659 7160 34704 7188
rect 34698 7148 34704 7160
rect 34756 7148 34762 7200
rect 1104 7098 58880 7120
rect 1104 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 8302 7098
rect 8354 7046 8366 7098
rect 8418 7046 8430 7098
rect 8482 7046 22622 7098
rect 22674 7046 22686 7098
rect 22738 7046 22750 7098
rect 22802 7046 22814 7098
rect 22866 7046 22878 7098
rect 22930 7046 37070 7098
rect 37122 7046 37134 7098
rect 37186 7046 37198 7098
rect 37250 7046 37262 7098
rect 37314 7046 37326 7098
rect 37378 7046 51518 7098
rect 51570 7046 51582 7098
rect 51634 7046 51646 7098
rect 51698 7046 51710 7098
rect 51762 7046 51774 7098
rect 51826 7046 58880 7098
rect 1104 7024 58880 7046
rect 21634 6984 21640 6996
rect 21595 6956 21640 6984
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 30466 6944 30472 6996
rect 30524 6984 30530 6996
rect 30561 6987 30619 6993
rect 30561 6984 30573 6987
rect 30524 6956 30573 6984
rect 30524 6944 30530 6956
rect 30561 6953 30573 6956
rect 30607 6953 30619 6987
rect 30561 6947 30619 6953
rect 31202 6944 31208 6996
rect 31260 6984 31266 6996
rect 31573 6987 31631 6993
rect 31573 6984 31585 6987
rect 31260 6956 31585 6984
rect 31260 6944 31266 6956
rect 31573 6953 31585 6956
rect 31619 6953 31631 6987
rect 31573 6947 31631 6953
rect 31665 6987 31723 6993
rect 31665 6953 31677 6987
rect 31711 6984 31723 6987
rect 31846 6984 31852 6996
rect 31711 6956 31852 6984
rect 31711 6953 31723 6956
rect 31665 6947 31723 6953
rect 31846 6944 31852 6956
rect 31904 6944 31910 6996
rect 33505 6987 33563 6993
rect 33505 6953 33517 6987
rect 33551 6984 33563 6987
rect 33778 6984 33784 6996
rect 33551 6956 33784 6984
rect 33551 6953 33563 6956
rect 33505 6947 33563 6953
rect 33778 6944 33784 6956
rect 33836 6944 33842 6996
rect 34698 6944 34704 6996
rect 34756 6984 34762 6996
rect 35602 6987 35660 6993
rect 35602 6984 35614 6987
rect 34756 6956 35614 6984
rect 34756 6944 34762 6956
rect 35602 6953 35614 6956
rect 35648 6953 35660 6987
rect 45094 6984 45100 6996
rect 45055 6956 45100 6984
rect 35602 6947 35660 6953
rect 45094 6944 45100 6956
rect 45152 6944 45158 6996
rect 45925 6987 45983 6993
rect 45925 6953 45937 6987
rect 45971 6984 45983 6987
rect 46382 6984 46388 6996
rect 45971 6956 46388 6984
rect 45971 6953 45983 6956
rect 45925 6947 45983 6953
rect 46382 6944 46388 6956
rect 46440 6944 46446 6996
rect 46474 6944 46480 6996
rect 46532 6984 46538 6996
rect 46532 6956 46577 6984
rect 46532 6944 46538 6956
rect 27982 6916 27988 6928
rect 27943 6888 27988 6916
rect 27982 6876 27988 6888
rect 28040 6876 28046 6928
rect 35066 6916 35072 6928
rect 33428 6888 35072 6916
rect 20349 6851 20407 6857
rect 20349 6817 20361 6851
rect 20395 6848 20407 6851
rect 20530 6848 20536 6860
rect 20395 6820 20536 6848
rect 20395 6817 20407 6820
rect 20349 6811 20407 6817
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 27614 6848 27620 6860
rect 27356 6820 27620 6848
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 19518 6780 19524 6792
rect 7984 6752 19524 6780
rect 7984 6740 7990 6752
rect 19518 6740 19524 6752
rect 19576 6780 19582 6792
rect 27356 6789 27384 6820
rect 27614 6808 27620 6820
rect 27672 6848 27678 6860
rect 27672 6820 28212 6848
rect 27672 6808 27678 6820
rect 20165 6783 20223 6789
rect 20165 6780 20177 6783
rect 19576 6752 20177 6780
rect 19576 6740 19582 6752
rect 20165 6749 20177 6752
rect 20211 6749 20223 6783
rect 20165 6743 20223 6749
rect 27341 6783 27399 6789
rect 27341 6749 27353 6783
rect 27387 6749 27399 6783
rect 27341 6743 27399 6749
rect 27525 6783 27583 6789
rect 27525 6749 27537 6783
rect 27571 6780 27583 6783
rect 27798 6780 27804 6792
rect 27571 6752 27804 6780
rect 27571 6749 27583 6752
rect 27525 6743 27583 6749
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 28184 6789 28212 6820
rect 29454 6808 29460 6860
rect 29512 6848 29518 6860
rect 31481 6851 31539 6857
rect 31481 6848 31493 6851
rect 29512 6820 31493 6848
rect 29512 6808 29518 6820
rect 31481 6817 31493 6820
rect 31527 6848 31539 6851
rect 31570 6848 31576 6860
rect 31527 6820 31576 6848
rect 31527 6817 31539 6820
rect 31481 6811 31539 6817
rect 31570 6808 31576 6820
rect 31628 6808 31634 6860
rect 32214 6848 32220 6860
rect 32175 6820 32220 6848
rect 32214 6808 32220 6820
rect 32272 6808 32278 6860
rect 28169 6783 28227 6789
rect 28169 6749 28181 6783
rect 28215 6749 28227 6783
rect 28169 6743 28227 6749
rect 29086 6740 29092 6792
rect 29144 6780 29150 6792
rect 29549 6783 29607 6789
rect 29549 6780 29561 6783
rect 29144 6752 29561 6780
rect 29144 6740 29150 6752
rect 29549 6749 29561 6752
rect 29595 6749 29607 6783
rect 29549 6743 29607 6749
rect 29733 6783 29791 6789
rect 29733 6749 29745 6783
rect 29779 6780 29791 6783
rect 30190 6780 30196 6792
rect 29779 6752 30196 6780
rect 29779 6749 29791 6752
rect 29733 6743 29791 6749
rect 30190 6740 30196 6752
rect 30248 6740 30254 6792
rect 30466 6780 30472 6792
rect 30427 6752 30472 6780
rect 30466 6740 30472 6752
rect 30524 6740 30530 6792
rect 30558 6740 30564 6792
rect 30616 6780 30622 6792
rect 30834 6780 30840 6792
rect 30616 6752 30661 6780
rect 30795 6752 30840 6780
rect 30616 6740 30622 6752
rect 30834 6740 30840 6752
rect 30892 6740 30898 6792
rect 33428 6789 33456 6888
rect 35066 6876 35072 6888
rect 35124 6876 35130 6928
rect 34238 6808 34244 6860
rect 34296 6848 34302 6860
rect 37093 6851 37151 6857
rect 37093 6848 37105 6851
rect 34296 6820 37105 6848
rect 34296 6808 34302 6820
rect 37093 6817 37105 6820
rect 37139 6817 37151 6851
rect 39022 6848 39028 6860
rect 38983 6820 39028 6848
rect 37093 6811 37151 6817
rect 39022 6808 39028 6820
rect 39080 6808 39086 6860
rect 39850 6808 39856 6860
rect 39908 6848 39914 6860
rect 40957 6851 41015 6857
rect 40957 6848 40969 6851
rect 39908 6820 40969 6848
rect 39908 6808 39914 6820
rect 40957 6817 40969 6820
rect 41003 6817 41015 6851
rect 40957 6811 41015 6817
rect 41800 6820 42656 6848
rect 31757 6783 31815 6789
rect 31757 6749 31769 6783
rect 31803 6780 31815 6783
rect 33413 6783 33471 6789
rect 33413 6780 33425 6783
rect 31803 6752 33425 6780
rect 31803 6749 31815 6752
rect 31757 6743 31815 6749
rect 33413 6749 33425 6752
rect 33459 6749 33471 6783
rect 33413 6743 33471 6749
rect 33597 6783 33655 6789
rect 33597 6749 33609 6783
rect 33643 6780 33655 6783
rect 34422 6780 34428 6792
rect 33643 6752 34428 6780
rect 33643 6749 33655 6752
rect 33597 6743 33655 6749
rect 28350 6712 28356 6724
rect 28263 6684 28356 6712
rect 28350 6672 28356 6684
rect 28408 6712 28414 6724
rect 31772 6712 31800 6743
rect 34422 6740 34428 6752
rect 34480 6740 34486 6792
rect 34514 6740 34520 6792
rect 34572 6780 34578 6792
rect 34701 6783 34759 6789
rect 34701 6780 34713 6783
rect 34572 6752 34713 6780
rect 34572 6740 34578 6752
rect 34701 6749 34713 6752
rect 34747 6749 34759 6783
rect 34701 6743 34759 6749
rect 35066 6740 35072 6792
rect 35124 6780 35130 6792
rect 35345 6783 35403 6789
rect 35345 6780 35357 6783
rect 35124 6752 35357 6780
rect 35124 6740 35130 6752
rect 35345 6749 35357 6752
rect 35391 6749 35403 6783
rect 35345 6743 35403 6749
rect 38197 6783 38255 6789
rect 38197 6749 38209 6783
rect 38243 6780 38255 6783
rect 38470 6780 38476 6792
rect 38243 6752 38476 6780
rect 38243 6749 38255 6752
rect 38197 6743 38255 6749
rect 38470 6740 38476 6752
rect 38528 6740 38534 6792
rect 38838 6740 38844 6792
rect 38896 6780 38902 6792
rect 38933 6783 38991 6789
rect 38933 6780 38945 6783
rect 38896 6752 38945 6780
rect 38896 6740 38902 6752
rect 38933 6749 38945 6752
rect 38979 6749 38991 6783
rect 39114 6780 39120 6792
rect 39075 6752 39120 6780
rect 38933 6743 38991 6749
rect 39114 6740 39120 6752
rect 39172 6740 39178 6792
rect 40402 6780 40408 6792
rect 40363 6752 40408 6780
rect 40402 6740 40408 6752
rect 40460 6740 40466 6792
rect 41800 6789 41828 6820
rect 42628 6789 42656 6820
rect 41785 6783 41843 6789
rect 41785 6749 41797 6783
rect 41831 6749 41843 6783
rect 41785 6743 41843 6749
rect 41969 6783 42027 6789
rect 41969 6749 41981 6783
rect 42015 6780 42027 6783
rect 42613 6783 42671 6789
rect 42015 6752 42472 6780
rect 42015 6749 42027 6752
rect 41969 6743 42027 6749
rect 38010 6712 38016 6724
rect 28408 6684 31800 6712
rect 36846 6684 38016 6712
rect 28408 6672 28414 6684
rect 38010 6672 38016 6684
rect 38068 6672 38074 6724
rect 40678 6672 40684 6724
rect 40736 6712 40742 6724
rect 41800 6712 41828 6743
rect 42444 6721 42472 6752
rect 42613 6749 42625 6783
rect 42659 6780 42671 6783
rect 44082 6780 44088 6792
rect 42659 6752 44088 6780
rect 42659 6749 42671 6752
rect 42613 6743 42671 6749
rect 44082 6740 44088 6752
rect 44140 6740 44146 6792
rect 45554 6740 45560 6792
rect 45612 6780 45618 6792
rect 45833 6783 45891 6789
rect 45833 6780 45845 6783
rect 45612 6752 45845 6780
rect 45612 6740 45618 6752
rect 45833 6749 45845 6752
rect 45879 6749 45891 6783
rect 45833 6743 45891 6749
rect 45922 6740 45928 6792
rect 45980 6780 45986 6792
rect 46017 6783 46075 6789
rect 46017 6780 46029 6783
rect 45980 6752 46029 6780
rect 45980 6740 45986 6752
rect 46017 6749 46029 6752
rect 46063 6780 46075 6783
rect 47029 6783 47087 6789
rect 47029 6780 47041 6783
rect 46063 6752 47041 6780
rect 46063 6749 46075 6752
rect 46017 6743 46075 6749
rect 47029 6749 47041 6752
rect 47075 6749 47087 6783
rect 47029 6743 47087 6749
rect 40736 6684 41828 6712
rect 42429 6715 42487 6721
rect 40736 6672 40742 6684
rect 42429 6681 42441 6715
rect 42475 6712 42487 6715
rect 43070 6712 43076 6724
rect 42475 6684 43076 6712
rect 42475 6681 42487 6684
rect 42429 6675 42487 6681
rect 43070 6672 43076 6684
rect 43128 6672 43134 6724
rect 43809 6715 43867 6721
rect 43809 6681 43821 6715
rect 43855 6712 43867 6715
rect 44726 6712 44732 6724
rect 43855 6684 44732 6712
rect 43855 6681 43867 6684
rect 43809 6675 43867 6681
rect 44726 6672 44732 6684
rect 44784 6672 44790 6724
rect 19702 6644 19708 6656
rect 19663 6616 19708 6644
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 27433 6647 27491 6653
rect 27433 6613 27445 6647
rect 27479 6644 27491 6647
rect 27706 6644 27712 6656
rect 27479 6616 27712 6644
rect 27479 6613 27491 6616
rect 27433 6607 27491 6613
rect 27706 6604 27712 6616
rect 27764 6604 27770 6656
rect 28258 6644 28264 6656
rect 28219 6616 28264 6644
rect 28258 6604 28264 6616
rect 28316 6604 28322 6656
rect 28537 6647 28595 6653
rect 28537 6613 28549 6647
rect 28583 6644 28595 6647
rect 29178 6644 29184 6656
rect 28583 6616 29184 6644
rect 28583 6613 28595 6616
rect 28537 6607 28595 6613
rect 29178 6604 29184 6616
rect 29236 6644 29242 6656
rect 29362 6644 29368 6656
rect 29236 6616 29368 6644
rect 29236 6604 29242 6616
rect 29362 6604 29368 6616
rect 29420 6604 29426 6656
rect 29730 6644 29736 6656
rect 29691 6616 29736 6644
rect 29730 6604 29736 6616
rect 29788 6604 29794 6656
rect 30650 6604 30656 6656
rect 30708 6644 30714 6656
rect 40313 6647 40371 6653
rect 30708 6616 30753 6644
rect 30708 6604 30714 6616
rect 40313 6613 40325 6647
rect 40359 6644 40371 6647
rect 40402 6644 40408 6656
rect 40359 6616 40408 6644
rect 40359 6613 40371 6616
rect 40313 6607 40371 6613
rect 40402 6604 40408 6616
rect 40460 6604 40466 6656
rect 41874 6644 41880 6656
rect 41835 6616 41880 6644
rect 41874 6604 41880 6616
rect 41932 6604 41938 6656
rect 42797 6647 42855 6653
rect 42797 6613 42809 6647
rect 42843 6644 42855 6647
rect 42886 6644 42892 6656
rect 42843 6616 42892 6644
rect 42843 6613 42855 6616
rect 42797 6607 42855 6613
rect 42886 6604 42892 6616
rect 42944 6604 42950 6656
rect 42978 6604 42984 6656
rect 43036 6644 43042 6656
rect 43717 6647 43775 6653
rect 43717 6644 43729 6647
rect 43036 6616 43729 6644
rect 43036 6604 43042 6616
rect 43717 6613 43729 6616
rect 43763 6613 43775 6647
rect 43717 6607 43775 6613
rect 1104 6554 58880 6576
rect 1104 6502 15398 6554
rect 15450 6502 15462 6554
rect 15514 6502 15526 6554
rect 15578 6502 15590 6554
rect 15642 6502 15654 6554
rect 15706 6502 29846 6554
rect 29898 6502 29910 6554
rect 29962 6502 29974 6554
rect 30026 6502 30038 6554
rect 30090 6502 30102 6554
rect 30154 6502 44294 6554
rect 44346 6502 44358 6554
rect 44410 6502 44422 6554
rect 44474 6502 44486 6554
rect 44538 6502 44550 6554
rect 44602 6502 58880 6554
rect 1104 6480 58880 6502
rect 19518 6440 19524 6452
rect 19479 6412 19524 6440
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 34422 6400 34428 6452
rect 34480 6440 34486 6452
rect 35069 6443 35127 6449
rect 35069 6440 35081 6443
rect 34480 6412 35081 6440
rect 34480 6400 34486 6412
rect 35069 6409 35081 6412
rect 35115 6409 35127 6443
rect 36722 6440 36728 6452
rect 36683 6412 36728 6440
rect 35069 6403 35127 6409
rect 36722 6400 36728 6412
rect 36780 6400 36786 6452
rect 41874 6400 41880 6452
rect 41932 6440 41938 6452
rect 42797 6443 42855 6449
rect 42797 6440 42809 6443
rect 41932 6412 42809 6440
rect 41932 6400 41938 6412
rect 42797 6409 42809 6412
rect 42843 6409 42855 6443
rect 42797 6403 42855 6409
rect 45649 6443 45707 6449
rect 45649 6409 45661 6443
rect 45695 6440 45707 6443
rect 45922 6440 45928 6452
rect 45695 6412 45928 6440
rect 45695 6409 45707 6412
rect 45649 6403 45707 6409
rect 45922 6400 45928 6412
rect 45980 6440 45986 6452
rect 46109 6443 46167 6449
rect 46109 6440 46121 6443
rect 45980 6412 46121 6440
rect 45980 6400 45986 6412
rect 46109 6409 46121 6412
rect 46155 6409 46167 6443
rect 46109 6403 46167 6409
rect 27157 6375 27215 6381
rect 27157 6341 27169 6375
rect 27203 6372 27215 6375
rect 27798 6372 27804 6384
rect 27203 6344 27804 6372
rect 27203 6341 27215 6344
rect 27157 6335 27215 6341
rect 27798 6332 27804 6344
rect 27856 6332 27862 6384
rect 28169 6375 28227 6381
rect 28169 6341 28181 6375
rect 28215 6372 28227 6375
rect 28258 6372 28264 6384
rect 28215 6344 28264 6372
rect 28215 6341 28227 6344
rect 28169 6335 28227 6341
rect 28258 6332 28264 6344
rect 28316 6372 28322 6384
rect 33594 6372 33600 6384
rect 28316 6344 31064 6372
rect 33555 6344 33600 6372
rect 28316 6332 28322 6344
rect 27709 6307 27767 6313
rect 27709 6273 27721 6307
rect 27755 6304 27767 6307
rect 28074 6304 28080 6316
rect 27755 6276 28080 6304
rect 27755 6273 27767 6276
rect 27709 6267 27767 6273
rect 28074 6264 28080 6276
rect 28132 6264 28138 6316
rect 29362 6304 29368 6316
rect 29275 6276 29368 6304
rect 29362 6264 29368 6276
rect 29420 6304 29426 6316
rect 30466 6304 30472 6316
rect 29420 6276 30472 6304
rect 29420 6264 29426 6276
rect 30466 6264 30472 6276
rect 30524 6264 30530 6316
rect 31036 6313 31064 6344
rect 33594 6332 33600 6344
rect 33652 6332 33658 6384
rect 35894 6372 35900 6384
rect 34822 6344 35900 6372
rect 35894 6332 35900 6344
rect 35952 6332 35958 6384
rect 36740 6372 36768 6400
rect 36740 6344 37780 6372
rect 31021 6307 31079 6313
rect 31021 6273 31033 6307
rect 31067 6304 31079 6307
rect 33226 6304 33232 6316
rect 31067 6276 33232 6304
rect 31067 6273 31079 6276
rect 31021 6267 31079 6273
rect 33226 6264 33232 6276
rect 33284 6264 33290 6316
rect 37752 6313 37780 6344
rect 38194 6332 38200 6384
rect 38252 6372 38258 6384
rect 41141 6375 41199 6381
rect 38252 6344 39068 6372
rect 38252 6332 38258 6344
rect 37737 6307 37795 6313
rect 37737 6273 37749 6307
rect 37783 6273 37795 6307
rect 37918 6304 37924 6316
rect 37879 6276 37924 6304
rect 37737 6267 37795 6273
rect 37918 6264 37924 6276
rect 37976 6264 37982 6316
rect 38746 6304 38752 6316
rect 38707 6276 38752 6304
rect 38746 6264 38752 6276
rect 38804 6264 38810 6316
rect 39040 6313 39068 6344
rect 41141 6341 41153 6375
rect 41187 6372 41199 6375
rect 41782 6372 41788 6384
rect 41187 6344 41788 6372
rect 41187 6341 41199 6344
rect 41141 6335 41199 6341
rect 41782 6332 41788 6344
rect 41840 6332 41846 6384
rect 44637 6375 44695 6381
rect 44637 6372 44649 6375
rect 42168 6344 44649 6372
rect 39025 6307 39083 6313
rect 39025 6273 39037 6307
rect 39071 6304 39083 6307
rect 39071 6276 39344 6304
rect 39071 6273 39083 6276
rect 39025 6267 39083 6273
rect 25958 6196 25964 6248
rect 26016 6236 26022 6248
rect 27065 6239 27123 6245
rect 27065 6236 27077 6239
rect 26016 6208 27077 6236
rect 26016 6196 26022 6208
rect 27065 6205 27077 6208
rect 27111 6205 27123 6239
rect 27065 6199 27123 6205
rect 29089 6239 29147 6245
rect 29089 6205 29101 6239
rect 29135 6236 29147 6239
rect 29454 6236 29460 6248
rect 29135 6208 29460 6236
rect 29135 6205 29147 6208
rect 29089 6199 29147 6205
rect 29454 6196 29460 6208
rect 29512 6196 29518 6248
rect 29730 6196 29736 6248
rect 29788 6236 29794 6248
rect 30929 6239 30987 6245
rect 30929 6236 30941 6239
rect 29788 6208 30941 6236
rect 29788 6196 29794 6208
rect 30929 6205 30941 6208
rect 30975 6205 30987 6239
rect 30929 6199 30987 6205
rect 32398 6196 32404 6248
rect 32456 6236 32462 6248
rect 33321 6239 33379 6245
rect 33321 6236 33333 6239
rect 32456 6208 33333 6236
rect 32456 6196 32462 6208
rect 33321 6205 33333 6208
rect 33367 6205 33379 6239
rect 33321 6199 33379 6205
rect 36630 6196 36636 6248
rect 36688 6236 36694 6248
rect 38841 6239 38899 6245
rect 38841 6236 38853 6239
rect 36688 6208 38853 6236
rect 36688 6196 36694 6208
rect 38841 6205 38853 6208
rect 38887 6205 38899 6239
rect 38841 6199 38899 6205
rect 27706 6128 27712 6180
rect 27764 6168 27770 6180
rect 28445 6171 28503 6177
rect 28445 6168 28457 6171
rect 27764 6140 28457 6168
rect 27764 6128 27770 6140
rect 28445 6137 28457 6140
rect 28491 6137 28503 6171
rect 28445 6131 28503 6137
rect 28629 6171 28687 6177
rect 28629 6137 28641 6171
rect 28675 6168 28687 6171
rect 29273 6171 29331 6177
rect 29273 6168 29285 6171
rect 28675 6140 29285 6168
rect 28675 6137 28687 6140
rect 28629 6131 28687 6137
rect 29273 6137 29285 6140
rect 29319 6137 29331 6171
rect 29273 6131 29331 6137
rect 31389 6171 31447 6177
rect 31389 6137 31401 6171
rect 31435 6168 31447 6171
rect 33226 6168 33232 6180
rect 31435 6140 33232 6168
rect 31435 6137 31447 6140
rect 31389 6131 31447 6137
rect 33226 6128 33232 6140
rect 33284 6128 33290 6180
rect 39209 6171 39267 6177
rect 39209 6168 39221 6171
rect 34624 6140 39221 6168
rect 28718 6060 28724 6112
rect 28776 6100 28782 6112
rect 29181 6103 29239 6109
rect 29181 6100 29193 6103
rect 28776 6072 29193 6100
rect 28776 6060 28782 6072
rect 29181 6069 29193 6072
rect 29227 6069 29239 6103
rect 29181 6063 29239 6069
rect 29917 6103 29975 6109
rect 29917 6069 29929 6103
rect 29963 6100 29975 6103
rect 30190 6100 30196 6112
rect 29963 6072 30196 6100
rect 29963 6069 29975 6072
rect 29917 6063 29975 6069
rect 30190 6060 30196 6072
rect 30248 6100 30254 6112
rect 32214 6100 32220 6112
rect 30248 6072 32220 6100
rect 30248 6060 30254 6072
rect 32214 6060 32220 6072
rect 32272 6060 32278 6112
rect 32582 6060 32588 6112
rect 32640 6100 32646 6112
rect 34624 6100 34652 6140
rect 39209 6137 39221 6140
rect 39255 6137 39267 6171
rect 39316 6168 39344 6276
rect 39850 6264 39856 6316
rect 39908 6304 39914 6316
rect 40221 6307 40279 6313
rect 40221 6304 40233 6307
rect 39908 6276 40233 6304
rect 39908 6264 39914 6276
rect 40221 6273 40233 6276
rect 40267 6273 40279 6307
rect 40221 6267 40279 6273
rect 41506 6264 41512 6316
rect 41564 6304 41570 6316
rect 41693 6307 41751 6313
rect 41693 6304 41705 6307
rect 41564 6276 41705 6304
rect 41564 6264 41570 6276
rect 41693 6273 41705 6276
rect 41739 6304 41751 6307
rect 42168 6304 42196 6344
rect 44637 6341 44649 6344
rect 44683 6341 44695 6375
rect 44637 6335 44695 6341
rect 41739 6276 42196 6304
rect 42705 6307 42763 6313
rect 41739 6273 41751 6276
rect 41693 6267 41751 6273
rect 42705 6273 42717 6307
rect 42751 6304 42763 6307
rect 42886 6304 42892 6316
rect 42751 6276 42892 6304
rect 42751 6273 42763 6276
rect 42705 6267 42763 6273
rect 42886 6264 42892 6276
rect 42944 6264 42950 6316
rect 42978 6264 42984 6316
rect 43036 6304 43042 6316
rect 43990 6304 43996 6316
rect 43036 6276 43081 6304
rect 43951 6276 43996 6304
rect 43036 6264 43042 6276
rect 43990 6264 43996 6276
rect 44048 6264 44054 6316
rect 40313 6239 40371 6245
rect 40313 6205 40325 6239
rect 40359 6236 40371 6239
rect 40678 6236 40684 6248
rect 40359 6208 40684 6236
rect 40359 6205 40371 6208
rect 40313 6199 40371 6205
rect 40678 6196 40684 6208
rect 40736 6236 40742 6248
rect 40957 6239 41015 6245
rect 40957 6236 40969 6239
rect 40736 6208 40969 6236
rect 40736 6196 40742 6208
rect 40957 6205 40969 6208
rect 41003 6205 41015 6239
rect 40957 6199 41015 6205
rect 43165 6239 43223 6245
rect 43165 6205 43177 6239
rect 43211 6236 43223 6239
rect 43901 6239 43959 6245
rect 43901 6236 43913 6239
rect 43211 6208 43913 6236
rect 43211 6205 43223 6208
rect 43165 6199 43223 6205
rect 43901 6205 43913 6208
rect 43947 6205 43959 6239
rect 43901 6199 43959 6205
rect 40586 6168 40592 6180
rect 39316 6140 40592 6168
rect 39209 6131 39267 6137
rect 40586 6128 40592 6140
rect 40644 6128 40650 6180
rect 43622 6168 43628 6180
rect 43583 6140 43628 6168
rect 43622 6128 43628 6140
rect 43680 6128 43686 6180
rect 32640 6072 34652 6100
rect 32640 6060 32646 6072
rect 37734 6060 37740 6112
rect 37792 6100 37798 6112
rect 37829 6103 37887 6109
rect 37829 6100 37841 6103
rect 37792 6072 37841 6100
rect 37792 6060 37798 6072
rect 37829 6069 37841 6072
rect 37875 6069 37887 6103
rect 39022 6100 39028 6112
rect 38983 6072 39028 6100
rect 37829 6063 37887 6069
rect 39022 6060 39028 6072
rect 39080 6060 39086 6112
rect 39853 6103 39911 6109
rect 39853 6069 39865 6103
rect 39899 6100 39911 6103
rect 40126 6100 40132 6112
rect 39899 6072 40132 6100
rect 39899 6069 39911 6072
rect 39853 6063 39911 6069
rect 40126 6060 40132 6072
rect 40184 6060 40190 6112
rect 41877 6103 41935 6109
rect 41877 6069 41889 6103
rect 41923 6100 41935 6103
rect 43070 6100 43076 6112
rect 41923 6072 43076 6100
rect 41923 6069 41935 6072
rect 41877 6063 41935 6069
rect 43070 6060 43076 6072
rect 43128 6100 43134 6112
rect 43530 6100 43536 6112
rect 43128 6072 43536 6100
rect 43128 6060 43134 6072
rect 43530 6060 43536 6072
rect 43588 6060 43594 6112
rect 1104 6010 58880 6032
rect 1104 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 8302 6010
rect 8354 5958 8366 6010
rect 8418 5958 8430 6010
rect 8482 5958 22622 6010
rect 22674 5958 22686 6010
rect 22738 5958 22750 6010
rect 22802 5958 22814 6010
rect 22866 5958 22878 6010
rect 22930 5958 37070 6010
rect 37122 5958 37134 6010
rect 37186 5958 37198 6010
rect 37250 5958 37262 6010
rect 37314 5958 37326 6010
rect 37378 5958 51518 6010
rect 51570 5958 51582 6010
rect 51634 5958 51646 6010
rect 51698 5958 51710 6010
rect 51762 5958 51774 6010
rect 51826 5958 58880 6010
rect 1104 5936 58880 5958
rect 25958 5896 25964 5908
rect 25919 5868 25964 5896
rect 25958 5856 25964 5868
rect 26016 5856 26022 5908
rect 27798 5856 27804 5908
rect 27856 5896 27862 5908
rect 27893 5899 27951 5905
rect 27893 5896 27905 5899
rect 27856 5868 27905 5896
rect 27856 5856 27862 5868
rect 27893 5865 27905 5868
rect 27939 5896 27951 5899
rect 28902 5896 28908 5908
rect 27939 5868 28908 5896
rect 27939 5865 27951 5868
rect 27893 5859 27951 5865
rect 28902 5856 28908 5868
rect 28960 5856 28966 5908
rect 32306 5856 32312 5908
rect 32364 5896 32370 5908
rect 32490 5896 32496 5908
rect 32364 5868 32496 5896
rect 32364 5856 32370 5868
rect 32490 5856 32496 5868
rect 32548 5896 32554 5908
rect 32548 5868 37412 5896
rect 32548 5856 32554 5868
rect 28997 5831 29055 5837
rect 28997 5797 29009 5831
rect 29043 5828 29055 5831
rect 29043 5800 32536 5828
rect 29043 5797 29055 5800
rect 28997 5791 29055 5797
rect 28718 5760 28724 5772
rect 28679 5732 28724 5760
rect 28718 5720 28724 5732
rect 28776 5720 28782 5772
rect 32398 5760 32404 5772
rect 30484 5732 31754 5760
rect 32359 5732 32404 5760
rect 25777 5695 25835 5701
rect 25777 5661 25789 5695
rect 25823 5692 25835 5695
rect 26234 5692 26240 5704
rect 25823 5664 26240 5692
rect 25823 5661 25835 5664
rect 25777 5655 25835 5661
rect 26234 5652 26240 5664
rect 26292 5652 26298 5704
rect 28626 5692 28632 5704
rect 28587 5664 28632 5692
rect 28626 5652 28632 5664
rect 28684 5652 28690 5704
rect 30484 5701 30512 5732
rect 30469 5695 30527 5701
rect 30469 5661 30481 5695
rect 30515 5661 30527 5695
rect 30742 5692 30748 5704
rect 30703 5664 30748 5692
rect 30469 5655 30527 5661
rect 30742 5652 30748 5664
rect 30800 5652 30806 5704
rect 30834 5652 30840 5704
rect 30892 5692 30898 5704
rect 31018 5692 31024 5704
rect 30892 5664 31024 5692
rect 30892 5652 30898 5664
rect 31018 5652 31024 5664
rect 31076 5692 31082 5704
rect 31389 5695 31447 5701
rect 31389 5692 31401 5695
rect 31076 5664 31401 5692
rect 31076 5652 31082 5664
rect 31389 5661 31401 5664
rect 31435 5661 31447 5695
rect 31726 5692 31754 5732
rect 32398 5720 32404 5732
rect 32456 5720 32462 5772
rect 32508 5760 32536 5800
rect 35066 5788 35072 5840
rect 35124 5828 35130 5840
rect 36357 5831 36415 5837
rect 36357 5828 36369 5831
rect 35124 5800 36369 5828
rect 35124 5788 35130 5800
rect 36357 5797 36369 5800
rect 36403 5797 36415 5831
rect 36357 5791 36415 5797
rect 32677 5763 32735 5769
rect 32677 5760 32689 5763
rect 32508 5732 32689 5760
rect 32677 5729 32689 5732
rect 32723 5729 32735 5763
rect 32677 5723 32735 5729
rect 32766 5720 32772 5772
rect 32824 5760 32830 5772
rect 36372 5760 36400 5791
rect 37277 5763 37335 5769
rect 37277 5760 37289 5763
rect 32824 5732 33916 5760
rect 36372 5732 37289 5760
rect 32824 5720 32830 5732
rect 32306 5692 32312 5704
rect 31726 5664 32312 5692
rect 31389 5655 31447 5661
rect 28644 5624 28672 5652
rect 31205 5627 31263 5633
rect 31205 5624 31217 5627
rect 28644 5596 31217 5624
rect 31205 5593 31217 5596
rect 31251 5593 31263 5627
rect 31205 5587 31263 5593
rect 29178 5516 29184 5568
rect 29236 5556 29242 5568
rect 30285 5559 30343 5565
rect 30285 5556 30297 5559
rect 29236 5528 30297 5556
rect 29236 5516 29242 5528
rect 30285 5525 30297 5528
rect 30331 5525 30343 5559
rect 30650 5556 30656 5568
rect 30611 5528 30656 5556
rect 30285 5519 30343 5525
rect 30650 5516 30656 5528
rect 30708 5516 30714 5568
rect 31404 5556 31432 5655
rect 32306 5652 32312 5664
rect 32364 5652 32370 5704
rect 33888 5692 33916 5732
rect 37277 5729 37289 5732
rect 37323 5729 37335 5763
rect 37384 5760 37412 5868
rect 37918 5856 37924 5908
rect 37976 5896 37982 5908
rect 39853 5899 39911 5905
rect 39853 5896 39865 5899
rect 37976 5868 39865 5896
rect 37976 5856 37982 5868
rect 39853 5865 39865 5868
rect 39899 5865 39911 5899
rect 39853 5859 39911 5865
rect 39022 5828 39028 5840
rect 38983 5800 39028 5828
rect 39022 5788 39028 5800
rect 39080 5788 39086 5840
rect 42978 5828 42984 5840
rect 39132 5800 42984 5828
rect 39132 5760 39160 5800
rect 37384 5732 39160 5760
rect 40497 5763 40555 5769
rect 37277 5723 37335 5729
rect 40497 5729 40509 5763
rect 40543 5760 40555 5763
rect 40586 5760 40592 5772
rect 40543 5732 40592 5760
rect 40543 5729 40555 5732
rect 40497 5723 40555 5729
rect 40586 5720 40592 5732
rect 40644 5720 40650 5772
rect 41325 5763 41383 5769
rect 41325 5729 41337 5763
rect 41371 5760 41383 5763
rect 42337 5763 42395 5769
rect 42337 5760 42349 5763
rect 41371 5732 42349 5760
rect 41371 5729 41383 5732
rect 41325 5723 41383 5729
rect 42337 5729 42349 5732
rect 42383 5729 42395 5763
rect 42337 5723 42395 5729
rect 36722 5692 36728 5704
rect 33888 5664 36728 5692
rect 36722 5652 36728 5664
rect 36780 5652 36786 5704
rect 40218 5652 40224 5704
rect 40276 5692 40282 5704
rect 40313 5695 40371 5701
rect 40313 5692 40325 5695
rect 40276 5664 40325 5692
rect 40276 5652 40282 5664
rect 40313 5661 40325 5664
rect 40359 5661 40371 5695
rect 40313 5655 40371 5661
rect 41233 5695 41291 5701
rect 41233 5661 41245 5695
rect 41279 5692 41291 5695
rect 41506 5692 41512 5704
rect 41279 5664 41512 5692
rect 41279 5661 41291 5664
rect 41233 5655 41291 5661
rect 41506 5652 41512 5664
rect 41564 5652 41570 5704
rect 42536 5701 42564 5800
rect 42978 5788 42984 5800
rect 43036 5788 43042 5840
rect 44085 5831 44143 5837
rect 44085 5797 44097 5831
rect 44131 5797 44143 5831
rect 44085 5791 44143 5797
rect 44100 5760 44128 5791
rect 42720 5732 44128 5760
rect 42720 5701 42748 5732
rect 42521 5695 42579 5701
rect 42521 5661 42533 5695
rect 42567 5661 42579 5695
rect 42521 5655 42579 5661
rect 42705 5695 42763 5701
rect 42705 5661 42717 5695
rect 42751 5661 42763 5695
rect 42705 5655 42763 5661
rect 42797 5695 42855 5701
rect 42797 5661 42809 5695
rect 42843 5692 42855 5695
rect 43625 5695 43683 5701
rect 43625 5692 43637 5695
rect 42843 5664 43637 5692
rect 42843 5661 42855 5664
rect 42797 5655 42855 5661
rect 43625 5661 43637 5664
rect 43671 5661 43683 5695
rect 44082 5692 44088 5704
rect 44043 5664 44088 5692
rect 43625 5655 43683 5661
rect 44082 5652 44088 5664
rect 44140 5652 44146 5704
rect 32214 5584 32220 5636
rect 32272 5624 32278 5636
rect 32766 5624 32772 5636
rect 32272 5596 32772 5624
rect 32272 5584 32278 5596
rect 32766 5584 32772 5596
rect 32824 5584 32830 5636
rect 34330 5624 34336 5636
rect 33902 5596 34336 5624
rect 34330 5584 34336 5596
rect 34388 5584 34394 5636
rect 35069 5627 35127 5633
rect 35069 5593 35081 5627
rect 35115 5593 35127 5627
rect 37550 5624 37556 5636
rect 37511 5596 37556 5624
rect 35069 5587 35127 5593
rect 34149 5559 34207 5565
rect 34149 5556 34161 5559
rect 31404 5528 34161 5556
rect 34149 5525 34161 5528
rect 34195 5525 34207 5559
rect 35084 5556 35112 5587
rect 37550 5584 37556 5596
rect 37608 5584 37614 5636
rect 38010 5584 38016 5636
rect 38068 5584 38074 5636
rect 42886 5584 42892 5636
rect 42944 5624 42950 5636
rect 43257 5627 43315 5633
rect 43257 5624 43269 5627
rect 42944 5596 43269 5624
rect 42944 5584 42950 5596
rect 43257 5593 43269 5596
rect 43303 5593 43315 5627
rect 43438 5624 43444 5636
rect 43399 5596 43444 5624
rect 43257 5587 43315 5593
rect 43438 5584 43444 5596
rect 43496 5584 43502 5636
rect 43530 5584 43536 5636
rect 43588 5624 43594 5636
rect 44177 5627 44235 5633
rect 44177 5624 44189 5627
rect 43588 5596 44189 5624
rect 43588 5584 43594 5596
rect 44177 5593 44189 5596
rect 44223 5593 44235 5627
rect 44177 5587 44235 5593
rect 44361 5627 44419 5633
rect 44361 5593 44373 5627
rect 44407 5593 44419 5627
rect 44361 5587 44419 5593
rect 38930 5556 38936 5568
rect 35084 5528 38936 5556
rect 34149 5519 34207 5525
rect 38930 5516 38936 5528
rect 38988 5516 38994 5568
rect 39942 5516 39948 5568
rect 40000 5556 40006 5568
rect 40221 5559 40279 5565
rect 40221 5556 40233 5559
rect 40000 5528 40233 5556
rect 40000 5516 40006 5528
rect 40221 5525 40233 5528
rect 40267 5525 40279 5559
rect 40221 5519 40279 5525
rect 41601 5559 41659 5565
rect 41601 5525 41613 5559
rect 41647 5556 41659 5559
rect 42702 5556 42708 5568
rect 41647 5528 42708 5556
rect 41647 5525 41659 5528
rect 41601 5519 41659 5525
rect 42702 5516 42708 5528
rect 42760 5516 42766 5568
rect 43456 5556 43484 5584
rect 43990 5556 43996 5568
rect 43456 5528 43996 5556
rect 43990 5516 43996 5528
rect 44048 5556 44054 5568
rect 44376 5556 44404 5587
rect 44048 5528 44404 5556
rect 44048 5516 44054 5528
rect 1104 5466 58880 5488
rect 1104 5414 15398 5466
rect 15450 5414 15462 5466
rect 15514 5414 15526 5466
rect 15578 5414 15590 5466
rect 15642 5414 15654 5466
rect 15706 5414 29846 5466
rect 29898 5414 29910 5466
rect 29962 5414 29974 5466
rect 30026 5414 30038 5466
rect 30090 5414 30102 5466
rect 30154 5414 44294 5466
rect 44346 5414 44358 5466
rect 44410 5414 44422 5466
rect 44474 5414 44486 5466
rect 44538 5414 44550 5466
rect 44602 5414 58880 5466
rect 1104 5392 58880 5414
rect 19702 5312 19708 5364
rect 19760 5352 19766 5364
rect 20625 5355 20683 5361
rect 20625 5352 20637 5355
rect 19760 5324 20637 5352
rect 19760 5312 19766 5324
rect 20625 5321 20637 5324
rect 20671 5321 20683 5355
rect 20625 5315 20683 5321
rect 21726 5312 21732 5364
rect 21784 5352 21790 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 21784 5324 21833 5352
rect 21784 5312 21790 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 26234 5352 26240 5364
rect 26195 5324 26240 5352
rect 21821 5315 21879 5321
rect 26234 5312 26240 5324
rect 26292 5312 26298 5364
rect 30650 5312 30656 5364
rect 30708 5352 30714 5364
rect 30929 5355 30987 5361
rect 30929 5352 30941 5355
rect 30708 5324 30941 5352
rect 30708 5312 30714 5324
rect 30929 5321 30941 5324
rect 30975 5321 30987 5355
rect 33318 5352 33324 5364
rect 33279 5324 33324 5352
rect 30929 5315 30987 5321
rect 33318 5312 33324 5324
rect 33376 5312 33382 5364
rect 37277 5355 37335 5361
rect 37277 5321 37289 5355
rect 37323 5352 37335 5355
rect 37550 5352 37556 5364
rect 37323 5324 37556 5352
rect 37323 5321 37335 5324
rect 37277 5315 37335 5321
rect 37550 5312 37556 5324
rect 37608 5312 37614 5364
rect 40034 5312 40040 5364
rect 40092 5352 40098 5364
rect 40310 5352 40316 5364
rect 40092 5324 40316 5352
rect 40092 5312 40098 5324
rect 40310 5312 40316 5324
rect 40368 5312 40374 5364
rect 41417 5355 41475 5361
rect 41417 5321 41429 5355
rect 41463 5352 41475 5355
rect 41506 5352 41512 5364
rect 41463 5324 41512 5352
rect 41463 5321 41475 5324
rect 41417 5315 41475 5321
rect 41506 5312 41512 5324
rect 41564 5352 41570 5364
rect 41564 5324 42932 5352
rect 41564 5312 41570 5324
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 21085 5219 21143 5225
rect 1719 5188 2268 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 2240 5089 2268 5188
rect 21085 5185 21097 5219
rect 21131 5216 21143 5219
rect 21744 5216 21772 5312
rect 30282 5244 30288 5296
rect 30340 5284 30346 5296
rect 30340 5256 32628 5284
rect 30340 5244 30346 5256
rect 32600 5228 32628 5256
rect 34330 5244 34336 5296
rect 34388 5284 34394 5296
rect 35713 5287 35771 5293
rect 35713 5284 35725 5287
rect 34388 5256 35725 5284
rect 34388 5244 34394 5256
rect 35713 5253 35725 5256
rect 35759 5284 35771 5287
rect 35802 5284 35808 5296
rect 35759 5256 35808 5284
rect 35759 5253 35771 5256
rect 35713 5247 35771 5253
rect 35802 5244 35808 5256
rect 35860 5244 35866 5296
rect 38930 5244 38936 5296
rect 38988 5284 38994 5296
rect 39025 5287 39083 5293
rect 39025 5284 39037 5287
rect 38988 5256 39037 5284
rect 38988 5244 38994 5256
rect 39025 5253 39037 5256
rect 39071 5253 39083 5287
rect 41598 5284 41604 5296
rect 41559 5256 41604 5284
rect 39025 5247 39083 5253
rect 41598 5244 41604 5256
rect 41656 5244 41662 5296
rect 41782 5284 41788 5296
rect 41743 5256 41788 5284
rect 41782 5244 41788 5256
rect 41840 5284 41846 5296
rect 41840 5256 42656 5284
rect 41840 5244 41846 5256
rect 25866 5216 25872 5228
rect 21131 5188 21772 5216
rect 25827 5188 25872 5216
rect 21131 5185 21143 5188
rect 21085 5179 21143 5185
rect 25866 5176 25872 5188
rect 25924 5176 25930 5228
rect 26053 5219 26111 5225
rect 26053 5216 26065 5219
rect 25976 5188 26065 5216
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5148 21327 5151
rect 25976 5148 26004 5188
rect 26053 5185 26065 5188
rect 26099 5216 26111 5219
rect 26970 5216 26976 5228
rect 26099 5188 26976 5216
rect 26099 5185 26111 5188
rect 26053 5179 26111 5185
rect 26970 5176 26976 5188
rect 27028 5176 27034 5228
rect 28721 5219 28779 5225
rect 28721 5185 28733 5219
rect 28767 5216 28779 5219
rect 28767 5188 29592 5216
rect 28767 5185 28779 5188
rect 28721 5179 28779 5185
rect 21315 5120 26004 5148
rect 28813 5151 28871 5157
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 28813 5117 28825 5151
rect 28859 5148 28871 5151
rect 29178 5148 29184 5160
rect 28859 5120 29184 5148
rect 28859 5117 28871 5120
rect 28813 5111 28871 5117
rect 29178 5108 29184 5120
rect 29236 5108 29242 5160
rect 29564 5157 29592 5188
rect 29638 5176 29644 5228
rect 29696 5216 29702 5228
rect 29825 5219 29883 5225
rect 29825 5216 29837 5219
rect 29696 5188 29837 5216
rect 29696 5176 29702 5188
rect 29825 5185 29837 5188
rect 29871 5185 29883 5219
rect 29825 5179 29883 5185
rect 30466 5176 30472 5228
rect 30524 5216 30530 5228
rect 30837 5219 30895 5225
rect 30837 5216 30849 5219
rect 30524 5188 30849 5216
rect 30524 5176 30530 5188
rect 30837 5185 30849 5188
rect 30883 5185 30895 5219
rect 31018 5216 31024 5228
rect 30979 5188 31024 5216
rect 30837 5179 30895 5185
rect 31018 5176 31024 5188
rect 31076 5176 31082 5228
rect 32306 5216 32312 5228
rect 32267 5188 32312 5216
rect 32306 5176 32312 5188
rect 32364 5176 32370 5228
rect 32490 5216 32496 5228
rect 32451 5188 32496 5216
rect 32490 5176 32496 5188
rect 32548 5176 32554 5228
rect 32582 5176 32588 5228
rect 32640 5216 32646 5228
rect 37642 5216 37648 5228
rect 32640 5188 32685 5216
rect 37603 5188 37648 5216
rect 32640 5176 32646 5188
rect 37642 5176 37648 5188
rect 37700 5176 37706 5228
rect 38102 5176 38108 5228
rect 38160 5216 38166 5228
rect 38565 5219 38623 5225
rect 38565 5216 38577 5219
rect 38160 5188 38577 5216
rect 38160 5176 38166 5188
rect 38565 5185 38577 5188
rect 38611 5216 38623 5219
rect 40218 5216 40224 5228
rect 38611 5188 40224 5216
rect 38611 5185 38623 5188
rect 38565 5179 38623 5185
rect 40218 5176 40224 5188
rect 40276 5216 40282 5228
rect 41233 5219 41291 5225
rect 41233 5216 41245 5219
rect 40276 5188 41245 5216
rect 40276 5176 40282 5188
rect 41233 5185 41245 5188
rect 41279 5185 41291 5219
rect 41506 5216 41512 5228
rect 41467 5188 41512 5216
rect 41233 5179 41291 5185
rect 41506 5176 41512 5188
rect 41564 5176 41570 5228
rect 42628 5225 42656 5256
rect 42904 5225 42932 5324
rect 42613 5219 42671 5225
rect 42613 5185 42625 5219
rect 42659 5185 42671 5219
rect 42613 5179 42671 5185
rect 42889 5219 42947 5225
rect 42889 5185 42901 5219
rect 42935 5216 42947 5219
rect 43070 5216 43076 5228
rect 42935 5188 43076 5216
rect 42935 5185 42947 5188
rect 42889 5179 42947 5185
rect 43070 5176 43076 5188
rect 43128 5176 43134 5228
rect 29549 5151 29607 5157
rect 29549 5117 29561 5151
rect 29595 5148 29607 5151
rect 30374 5148 30380 5160
rect 29595 5120 30380 5148
rect 29595 5117 29607 5120
rect 29549 5111 29607 5117
rect 30374 5108 30380 5120
rect 30432 5148 30438 5160
rect 30558 5148 30564 5160
rect 30432 5120 30564 5148
rect 30432 5108 30438 5120
rect 30558 5108 30564 5120
rect 30616 5108 30622 5160
rect 31478 5108 31484 5160
rect 31536 5148 31542 5160
rect 32030 5148 32036 5160
rect 31536 5120 32036 5148
rect 31536 5108 31542 5120
rect 32030 5108 32036 5120
rect 32088 5148 32094 5160
rect 32088 5120 33180 5148
rect 32088 5108 32094 5120
rect 2225 5083 2283 5089
rect 2225 5049 2237 5083
rect 2271 5080 2283 5083
rect 24762 5080 24768 5092
rect 2271 5052 24768 5080
rect 2271 5049 2283 5052
rect 2225 5043 2283 5049
rect 24762 5040 24768 5052
rect 24820 5040 24826 5092
rect 29089 5083 29147 5089
rect 29089 5049 29101 5083
rect 29135 5080 29147 5083
rect 33042 5080 33048 5092
rect 29135 5052 33048 5080
rect 29135 5049 29147 5052
rect 29089 5043 29147 5049
rect 33042 5040 33048 5052
rect 33100 5040 33106 5092
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 24854 4972 24860 5024
rect 24912 5012 24918 5024
rect 25041 5015 25099 5021
rect 25041 5012 25053 5015
rect 24912 4984 25053 5012
rect 24912 4972 24918 4984
rect 25041 4981 25053 4984
rect 25087 4981 25099 5015
rect 32122 5012 32128 5024
rect 32083 4984 32128 5012
rect 25041 4975 25099 4981
rect 32122 4972 32128 4984
rect 32180 4972 32186 5024
rect 33152 5012 33180 5120
rect 33226 5108 33232 5160
rect 33284 5148 33290 5160
rect 34793 5151 34851 5157
rect 34793 5148 34805 5151
rect 33284 5120 34805 5148
rect 33284 5108 33290 5120
rect 34793 5117 34805 5120
rect 34839 5117 34851 5151
rect 35066 5148 35072 5160
rect 35027 5120 35072 5148
rect 34793 5111 34851 5117
rect 35066 5108 35072 5120
rect 35124 5108 35130 5160
rect 37734 5148 37740 5160
rect 37695 5120 37740 5148
rect 37734 5108 37740 5120
rect 37792 5108 37798 5160
rect 38286 5148 38292 5160
rect 38247 5120 38292 5148
rect 38286 5108 38292 5120
rect 38344 5108 38350 5160
rect 41524 5148 41552 5176
rect 42705 5151 42763 5157
rect 42705 5148 42717 5151
rect 41524 5120 42717 5148
rect 42705 5117 42717 5120
rect 42751 5148 42763 5151
rect 43438 5148 43444 5160
rect 42751 5120 43444 5148
rect 42751 5117 42763 5120
rect 42705 5111 42763 5117
rect 43438 5108 43444 5120
rect 43496 5108 43502 5160
rect 35250 5040 35256 5092
rect 35308 5080 35314 5092
rect 35529 5083 35587 5089
rect 35529 5080 35541 5083
rect 35308 5052 35541 5080
rect 35308 5040 35314 5052
rect 35529 5049 35541 5052
rect 35575 5049 35587 5083
rect 35529 5043 35587 5049
rect 39850 5040 39856 5092
rect 39908 5080 39914 5092
rect 39908 5052 41414 5080
rect 39908 5040 39914 5052
rect 36630 5012 36636 5024
rect 33152 4984 36636 5012
rect 36630 4972 36636 4984
rect 36688 4972 36694 5024
rect 37550 4972 37556 5024
rect 37608 5012 37614 5024
rect 38381 5015 38439 5021
rect 38381 5012 38393 5015
rect 37608 4984 38393 5012
rect 37608 4972 37614 4984
rect 38381 4981 38393 4984
rect 38427 4981 38439 5015
rect 38381 4975 38439 4981
rect 38473 5015 38531 5021
rect 38473 4981 38485 5015
rect 38519 5012 38531 5015
rect 39942 5012 39948 5024
rect 38519 4984 39948 5012
rect 38519 4981 38531 4984
rect 38473 4975 38531 4981
rect 39942 4972 39948 4984
rect 40000 4972 40006 5024
rect 41386 5012 41414 5052
rect 42429 5015 42487 5021
rect 42429 5012 42441 5015
rect 41386 4984 42441 5012
rect 42429 4981 42441 4984
rect 42475 4981 42487 5015
rect 42429 4975 42487 4981
rect 42889 5015 42947 5021
rect 42889 4981 42901 5015
rect 42935 5012 42947 5015
rect 43530 5012 43536 5024
rect 42935 4984 43536 5012
rect 42935 4981 42947 4984
rect 42889 4975 42947 4981
rect 43530 4972 43536 4984
rect 43588 4972 43594 5024
rect 1104 4922 58880 4944
rect 1104 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 8302 4922
rect 8354 4870 8366 4922
rect 8418 4870 8430 4922
rect 8482 4870 22622 4922
rect 22674 4870 22686 4922
rect 22738 4870 22750 4922
rect 22802 4870 22814 4922
rect 22866 4870 22878 4922
rect 22930 4870 37070 4922
rect 37122 4870 37134 4922
rect 37186 4870 37198 4922
rect 37250 4870 37262 4922
rect 37314 4870 37326 4922
rect 37378 4870 51518 4922
rect 51570 4870 51582 4922
rect 51634 4870 51646 4922
rect 51698 4870 51710 4922
rect 51762 4870 51774 4922
rect 51826 4870 58880 4922
rect 1104 4848 58880 4870
rect 24762 4808 24768 4820
rect 24723 4780 24768 4808
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 25866 4808 25872 4820
rect 25827 4780 25872 4808
rect 25866 4768 25872 4780
rect 25924 4768 25930 4820
rect 31021 4811 31079 4817
rect 31021 4808 31033 4811
rect 30668 4780 31033 4808
rect 25777 4743 25835 4749
rect 25777 4709 25789 4743
rect 25823 4740 25835 4743
rect 26326 4740 26332 4752
rect 25823 4712 26332 4740
rect 25823 4709 25835 4712
rect 25777 4703 25835 4709
rect 26326 4700 26332 4712
rect 26384 4700 26390 4752
rect 26605 4743 26663 4749
rect 26605 4709 26617 4743
rect 26651 4709 26663 4743
rect 26605 4703 26663 4709
rect 26620 4672 26648 4703
rect 27249 4675 27307 4681
rect 27249 4672 27261 4675
rect 25424 4644 27261 4672
rect 24854 4604 24860 4616
rect 24815 4576 24860 4604
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 25424 4548 25452 4644
rect 27249 4641 27261 4644
rect 27295 4641 27307 4675
rect 27249 4635 27307 4641
rect 28721 4675 28779 4681
rect 28721 4641 28733 4675
rect 28767 4672 28779 4675
rect 29638 4672 29644 4684
rect 28767 4644 29644 4672
rect 28767 4641 28779 4644
rect 28721 4635 28779 4641
rect 29638 4632 29644 4644
rect 29696 4632 29702 4684
rect 28997 4607 29055 4613
rect 28997 4573 29009 4607
rect 29043 4604 29055 4607
rect 29178 4604 29184 4616
rect 29043 4576 29184 4604
rect 29043 4573 29055 4576
rect 28997 4567 29055 4573
rect 29178 4564 29184 4576
rect 29236 4564 29242 4616
rect 25406 4536 25412 4548
rect 25367 4508 25412 4536
rect 25406 4496 25412 4508
rect 25464 4496 25470 4548
rect 26326 4536 26332 4548
rect 26287 4508 26332 4536
rect 26326 4496 26332 4508
rect 26384 4496 26390 4548
rect 30668 4536 30696 4780
rect 31021 4777 31033 4780
rect 31067 4777 31079 4811
rect 31021 4771 31079 4777
rect 31941 4811 31999 4817
rect 31941 4777 31953 4811
rect 31987 4808 31999 4811
rect 32490 4808 32496 4820
rect 31987 4780 32496 4808
rect 31987 4777 31999 4780
rect 31941 4771 31999 4777
rect 32490 4768 32496 4780
rect 32548 4768 32554 4820
rect 33134 4768 33140 4820
rect 33192 4808 33198 4820
rect 33965 4811 34023 4817
rect 33965 4808 33977 4811
rect 33192 4780 33977 4808
rect 33192 4768 33198 4780
rect 33965 4777 33977 4780
rect 34011 4777 34023 4811
rect 33965 4771 34023 4777
rect 37553 4811 37611 4817
rect 37553 4777 37565 4811
rect 37599 4808 37611 4811
rect 37642 4808 37648 4820
rect 37599 4780 37648 4808
rect 37599 4777 37611 4780
rect 37553 4771 37611 4777
rect 37642 4768 37648 4780
rect 37700 4808 37706 4820
rect 39942 4808 39948 4820
rect 37700 4780 38608 4808
rect 39903 4780 39948 4808
rect 37700 4768 37706 4780
rect 33321 4743 33379 4749
rect 33321 4740 33333 4743
rect 30852 4712 33333 4740
rect 30852 4681 30880 4712
rect 33321 4709 33333 4712
rect 33367 4709 33379 4743
rect 33321 4703 33379 4709
rect 33413 4743 33471 4749
rect 33413 4709 33425 4743
rect 33459 4740 33471 4743
rect 38473 4743 38531 4749
rect 38473 4740 38485 4743
rect 33459 4712 38485 4740
rect 33459 4709 33471 4712
rect 33413 4703 33471 4709
rect 38473 4709 38485 4712
rect 38519 4709 38531 4743
rect 38473 4703 38531 4709
rect 30837 4675 30895 4681
rect 30837 4641 30849 4675
rect 30883 4641 30895 4675
rect 30837 4635 30895 4641
rect 31386 4632 31392 4684
rect 31444 4672 31450 4684
rect 31444 4644 31754 4672
rect 31444 4632 31450 4644
rect 30745 4607 30803 4613
rect 30745 4573 30757 4607
rect 30791 4604 30803 4607
rect 31478 4604 31484 4616
rect 30791 4576 31484 4604
rect 30791 4573 30803 4576
rect 30745 4567 30803 4573
rect 31478 4564 31484 4576
rect 31536 4564 31542 4616
rect 31726 4604 31754 4644
rect 31864 4644 32168 4672
rect 31864 4613 31892 4644
rect 31849 4607 31907 4613
rect 31849 4604 31861 4607
rect 31726 4576 31861 4604
rect 31849 4573 31861 4576
rect 31895 4573 31907 4607
rect 32030 4604 32036 4616
rect 31991 4576 32036 4604
rect 31849 4567 31907 4573
rect 32030 4564 32036 4576
rect 32088 4564 32094 4616
rect 32140 4604 32168 4644
rect 33134 4632 33140 4684
rect 33192 4672 33198 4684
rect 33229 4675 33287 4681
rect 33229 4672 33241 4675
rect 33192 4644 33241 4672
rect 33192 4632 33198 4644
rect 33229 4641 33241 4644
rect 33275 4641 33287 4675
rect 38194 4672 38200 4684
rect 38155 4644 38200 4672
rect 33229 4635 33287 4641
rect 38194 4632 38200 4644
rect 38252 4632 38258 4684
rect 38381 4675 38439 4681
rect 38381 4641 38393 4675
rect 38427 4672 38439 4675
rect 38580 4672 38608 4780
rect 39942 4768 39948 4780
rect 40000 4768 40006 4820
rect 41506 4768 41512 4820
rect 41564 4808 41570 4820
rect 41693 4811 41751 4817
rect 41693 4808 41705 4811
rect 41564 4780 41705 4808
rect 41564 4768 41570 4780
rect 41693 4777 41705 4780
rect 41739 4777 41751 4811
rect 41693 4771 41751 4777
rect 41141 4743 41199 4749
rect 41141 4709 41153 4743
rect 41187 4740 41199 4743
rect 41598 4740 41604 4752
rect 41187 4712 41604 4740
rect 41187 4709 41199 4712
rect 41141 4703 41199 4709
rect 41598 4700 41604 4712
rect 41656 4700 41662 4752
rect 39022 4672 39028 4684
rect 38427 4644 39028 4672
rect 38427 4641 38439 4644
rect 38381 4635 38439 4641
rect 39022 4632 39028 4644
rect 39080 4632 39086 4684
rect 42426 4632 42432 4684
rect 42484 4672 42490 4684
rect 43441 4675 43499 4681
rect 43441 4672 43453 4675
rect 42484 4644 43453 4672
rect 42484 4632 42490 4644
rect 43441 4641 43453 4644
rect 43487 4641 43499 4675
rect 43441 4635 43499 4641
rect 33505 4607 33563 4613
rect 33505 4604 33517 4607
rect 32140 4576 33517 4604
rect 33505 4573 33517 4576
rect 33551 4604 33563 4607
rect 38102 4604 38108 4616
rect 33551 4576 37412 4604
rect 33551 4573 33563 4576
rect 33505 4567 33563 4573
rect 31754 4536 31760 4548
rect 28290 4508 29776 4536
rect 30668 4508 31760 4536
rect 26789 4471 26847 4477
rect 26789 4437 26801 4471
rect 26835 4468 26847 4471
rect 27154 4468 27160 4480
rect 26835 4440 27160 4468
rect 26835 4437 26847 4440
rect 26789 4431 26847 4437
rect 27154 4428 27160 4440
rect 27212 4428 27218 4480
rect 27246 4428 27252 4480
rect 27304 4468 27310 4480
rect 28368 4468 28396 4508
rect 29638 4468 29644 4480
rect 27304 4440 28396 4468
rect 29599 4440 29644 4468
rect 27304 4428 27310 4440
rect 29638 4428 29644 4440
rect 29696 4428 29702 4480
rect 29748 4468 29776 4508
rect 31754 4496 31760 4508
rect 31812 4496 31818 4548
rect 35069 4539 35127 4545
rect 35069 4536 35081 4539
rect 31864 4508 35081 4536
rect 31864 4468 31892 4508
rect 35069 4505 35081 4508
rect 35115 4505 35127 4539
rect 35250 4536 35256 4548
rect 35211 4508 35256 4536
rect 35069 4499 35127 4505
rect 35250 4496 35256 4508
rect 35308 4496 35314 4548
rect 37384 4477 37412 4576
rect 37660 4576 38108 4604
rect 37537 4539 37595 4545
rect 37537 4505 37549 4539
rect 37583 4536 37595 4539
rect 37660 4536 37688 4576
rect 38102 4564 38108 4576
rect 38160 4564 38166 4616
rect 37583 4508 37688 4536
rect 37583 4505 37595 4508
rect 37537 4499 37595 4505
rect 37734 4496 37740 4548
rect 37792 4536 37798 4548
rect 38212 4536 38240 4632
rect 38473 4607 38531 4613
rect 38473 4573 38485 4607
rect 38519 4604 38531 4607
rect 38746 4604 38752 4616
rect 38519 4576 38752 4604
rect 38519 4573 38531 4576
rect 38473 4567 38531 4573
rect 38746 4564 38752 4576
rect 38804 4604 38810 4616
rect 39850 4604 39856 4616
rect 38804 4576 39856 4604
rect 38804 4564 38810 4576
rect 39850 4564 39856 4576
rect 39908 4604 39914 4616
rect 40037 4607 40095 4613
rect 40037 4604 40049 4607
rect 39908 4576 40049 4604
rect 39908 4564 39914 4576
rect 40037 4573 40049 4576
rect 40083 4573 40095 4607
rect 40037 4567 40095 4573
rect 37792 4508 38240 4536
rect 37792 4496 37798 4508
rect 41322 4496 41328 4548
rect 41380 4536 41386 4548
rect 43165 4539 43223 4545
rect 41380 4508 41998 4536
rect 41380 4496 41386 4508
rect 43165 4505 43177 4539
rect 43211 4536 43223 4539
rect 43622 4536 43628 4548
rect 43211 4508 43628 4536
rect 43211 4505 43223 4508
rect 43165 4499 43223 4505
rect 43622 4496 43628 4508
rect 43680 4496 43686 4548
rect 29748 4440 31892 4468
rect 37369 4471 37427 4477
rect 37369 4437 37381 4471
rect 37415 4437 37427 4471
rect 37369 4431 37427 4437
rect 1104 4378 58880 4400
rect 1104 4326 15398 4378
rect 15450 4326 15462 4378
rect 15514 4326 15526 4378
rect 15578 4326 15590 4378
rect 15642 4326 15654 4378
rect 15706 4326 29846 4378
rect 29898 4326 29910 4378
rect 29962 4326 29974 4378
rect 30026 4326 30038 4378
rect 30090 4326 30102 4378
rect 30154 4326 44294 4378
rect 44346 4326 44358 4378
rect 44410 4326 44422 4378
rect 44474 4326 44486 4378
rect 44538 4326 44550 4378
rect 44602 4326 58880 4378
rect 1104 4304 58880 4326
rect 26970 4264 26976 4276
rect 26931 4236 26976 4264
rect 26970 4224 26976 4236
rect 27028 4224 27034 4276
rect 31754 4224 31760 4276
rect 31812 4264 31818 4276
rect 34422 4264 34428 4276
rect 31812 4236 34428 4264
rect 31812 4224 31818 4236
rect 34422 4224 34428 4236
rect 34480 4224 34486 4276
rect 35250 4264 35256 4276
rect 34808 4236 35256 4264
rect 27246 4196 27252 4208
rect 24150 4168 27252 4196
rect 27246 4156 27252 4168
rect 27304 4156 27310 4208
rect 34808 4196 34836 4236
rect 35250 4224 35256 4236
rect 35308 4224 35314 4276
rect 40586 4264 40592 4276
rect 40547 4236 40592 4264
rect 40586 4224 40592 4236
rect 40644 4224 40650 4276
rect 34178 4168 34836 4196
rect 35268 4196 35296 4224
rect 39117 4199 39175 4205
rect 39117 4196 39129 4199
rect 35268 4168 35650 4196
rect 38856 4168 39129 4196
rect 13630 4088 13636 4140
rect 13688 4128 13694 4140
rect 14274 4128 14280 4140
rect 13688 4100 14280 4128
rect 13688 4088 13694 4100
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 27154 4128 27160 4140
rect 27115 4100 27160 4128
rect 27154 4088 27160 4100
rect 27212 4088 27218 4140
rect 31021 4131 31079 4137
rect 31021 4097 31033 4131
rect 31067 4097 31079 4131
rect 32122 4128 32128 4140
rect 31021 4091 31079 4097
rect 31128 4100 32128 4128
rect 24581 4063 24639 4069
rect 24581 4029 24593 4063
rect 24627 4060 24639 4063
rect 24857 4063 24915 4069
rect 24627 4032 24808 4060
rect 24627 4029 24639 4032
rect 24581 4023 24639 4029
rect 24780 3992 24808 4032
rect 24857 4029 24869 4063
rect 24903 4060 24915 4063
rect 25314 4060 25320 4072
rect 24903 4032 25320 4060
rect 24903 4029 24915 4032
rect 24857 4023 24915 4029
rect 25314 4020 25320 4032
rect 25372 4020 25378 4072
rect 25406 3992 25412 4004
rect 24780 3964 25412 3992
rect 25406 3952 25412 3964
rect 25464 3952 25470 4004
rect 23106 3924 23112 3936
rect 23067 3896 23112 3924
rect 23106 3884 23112 3896
rect 23164 3884 23170 3936
rect 25314 3924 25320 3936
rect 25275 3896 25320 3924
rect 25314 3884 25320 3896
rect 25372 3884 25378 3936
rect 29178 3924 29184 3936
rect 29139 3896 29184 3924
rect 29178 3884 29184 3896
rect 29236 3884 29242 3936
rect 31036 3924 31064 4091
rect 31128 4069 31156 4100
rect 32122 4088 32128 4100
rect 32180 4088 32186 4140
rect 32398 4088 32404 4140
rect 32456 4128 32462 4140
rect 32677 4131 32735 4137
rect 32677 4128 32689 4131
rect 32456 4100 32689 4128
rect 32456 4088 32462 4100
rect 32677 4097 32689 4100
rect 32723 4097 32735 4131
rect 32677 4091 32735 4097
rect 37461 4131 37519 4137
rect 37461 4097 37473 4131
rect 37507 4128 37519 4131
rect 37734 4128 37740 4140
rect 37507 4100 37740 4128
rect 37507 4097 37519 4100
rect 37461 4091 37519 4097
rect 37734 4088 37740 4100
rect 37792 4088 37798 4140
rect 38856 4128 38884 4168
rect 39117 4165 39129 4168
rect 39163 4165 39175 4199
rect 40402 4196 40408 4208
rect 40342 4168 40408 4196
rect 39117 4159 39175 4165
rect 40402 4156 40408 4168
rect 40460 4196 40466 4208
rect 41322 4196 41328 4208
rect 40460 4168 41328 4196
rect 40460 4156 40466 4168
rect 41322 4156 41328 4168
rect 41380 4196 41386 4208
rect 41380 4168 43194 4196
rect 41380 4156 41386 4168
rect 42426 4128 42432 4140
rect 38396 4100 38884 4128
rect 41386 4100 42432 4128
rect 31113 4063 31171 4069
rect 31113 4029 31125 4063
rect 31159 4029 31171 4063
rect 32953 4063 33011 4069
rect 32953 4060 32965 4063
rect 31113 4023 31171 4029
rect 31726 4032 32965 4060
rect 31389 3995 31447 4001
rect 31389 3961 31401 3995
rect 31435 3992 31447 3995
rect 31726 3992 31754 4032
rect 32953 4029 32965 4032
rect 32999 4029 33011 4063
rect 34882 4060 34888 4072
rect 34843 4032 34888 4060
rect 32953 4023 33011 4029
rect 34882 4020 34888 4032
rect 34940 4020 34946 4072
rect 35161 4063 35219 4069
rect 35161 4060 35173 4063
rect 34992 4032 35173 4060
rect 31435 3964 31754 3992
rect 31435 3961 31447 3964
rect 31389 3955 31447 3961
rect 34514 3952 34520 4004
rect 34572 3992 34578 4004
rect 34992 3992 35020 4032
rect 35161 4029 35173 4032
rect 35207 4029 35219 4063
rect 36630 4060 36636 4072
rect 36591 4032 36636 4060
rect 35161 4023 35219 4029
rect 36630 4020 36636 4032
rect 36688 4020 36694 4072
rect 37550 4060 37556 4072
rect 37511 4032 37556 4060
rect 37550 4020 37556 4032
rect 37608 4020 37614 4072
rect 34572 3964 35020 3992
rect 37829 3995 37887 4001
rect 34572 3952 34578 3964
rect 37829 3961 37841 3995
rect 37875 3992 37887 3995
rect 38396 3992 38424 4100
rect 38841 4063 38899 4069
rect 38841 4029 38853 4063
rect 38887 4060 38899 4063
rect 40310 4060 40316 4072
rect 38887 4032 40316 4060
rect 38887 4029 38899 4032
rect 38841 4023 38899 4029
rect 40310 4020 40316 4032
rect 40368 4060 40374 4072
rect 41386 4060 41414 4100
rect 42426 4088 42432 4100
rect 42484 4088 42490 4140
rect 48682 4128 48688 4140
rect 48643 4100 48688 4128
rect 48682 4088 48688 4100
rect 48740 4128 48746 4140
rect 49329 4131 49387 4137
rect 49329 4128 49341 4131
rect 48740 4100 49341 4128
rect 48740 4088 48746 4100
rect 49329 4097 49341 4100
rect 49375 4097 49387 4131
rect 49329 4091 49387 4097
rect 42702 4060 42708 4072
rect 40368 4032 41414 4060
rect 42663 4032 42708 4060
rect 40368 4020 40374 4032
rect 42702 4020 42708 4032
rect 42760 4020 42766 4072
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 44177 4063 44235 4069
rect 44177 4060 44189 4063
rect 43128 4032 44189 4060
rect 43128 4020 43134 4032
rect 44177 4029 44189 4032
rect 44223 4029 44235 4063
rect 44177 4023 44235 4029
rect 37875 3964 38424 3992
rect 37875 3961 37887 3964
rect 37829 3955 37887 3961
rect 31938 3924 31944 3936
rect 31036 3896 31944 3924
rect 31938 3884 31944 3896
rect 31996 3924 32002 3936
rect 32582 3924 32588 3936
rect 31996 3896 32588 3924
rect 31996 3884 32002 3896
rect 32582 3884 32588 3896
rect 32640 3884 32646 3936
rect 34422 3884 34428 3936
rect 34480 3924 34486 3936
rect 48866 3924 48872 3936
rect 34480 3896 34525 3924
rect 48827 3896 48872 3924
rect 34480 3884 34486 3896
rect 48866 3884 48872 3896
rect 48924 3884 48930 3936
rect 1104 3834 58880 3856
rect 1104 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 8302 3834
rect 8354 3782 8366 3834
rect 8418 3782 8430 3834
rect 8482 3782 22622 3834
rect 22674 3782 22686 3834
rect 22738 3782 22750 3834
rect 22802 3782 22814 3834
rect 22866 3782 22878 3834
rect 22930 3782 37070 3834
rect 37122 3782 37134 3834
rect 37186 3782 37198 3834
rect 37250 3782 37262 3834
rect 37314 3782 37326 3834
rect 37378 3782 51518 3834
rect 51570 3782 51582 3834
rect 51634 3782 51646 3834
rect 51698 3782 51710 3834
rect 51762 3782 51774 3834
rect 51826 3782 58880 3834
rect 1104 3760 58880 3782
rect 26326 3680 26332 3732
rect 26384 3720 26390 3732
rect 27157 3723 27215 3729
rect 27157 3720 27169 3723
rect 26384 3692 27169 3720
rect 26384 3680 26390 3692
rect 27157 3689 27169 3692
rect 27203 3689 27215 3723
rect 27157 3683 27215 3689
rect 27709 3723 27767 3729
rect 27709 3689 27721 3723
rect 27755 3720 27767 3723
rect 29178 3720 29184 3732
rect 27755 3692 29184 3720
rect 27755 3689 27767 3692
rect 27709 3683 27767 3689
rect 23106 3544 23112 3596
rect 23164 3584 23170 3596
rect 25685 3587 25743 3593
rect 25685 3584 25697 3587
rect 23164 3556 25697 3584
rect 23164 3544 23170 3556
rect 25685 3553 25697 3556
rect 25731 3553 25743 3587
rect 25685 3547 25743 3553
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 25409 3519 25467 3525
rect 25409 3516 25421 3519
rect 25372 3488 25421 3516
rect 25372 3476 25378 3488
rect 25409 3485 25421 3488
rect 25455 3485 25467 3519
rect 25409 3479 25467 3485
rect 25424 3380 25452 3479
rect 27246 3448 27252 3460
rect 26910 3420 27252 3448
rect 27246 3408 27252 3420
rect 27304 3408 27310 3460
rect 27724 3380 27752 3683
rect 29178 3680 29184 3692
rect 29236 3680 29242 3732
rect 32582 3680 32588 3732
rect 32640 3720 32646 3732
rect 34422 3720 34428 3732
rect 32640 3692 34428 3720
rect 32640 3680 32646 3692
rect 34422 3680 34428 3692
rect 34480 3680 34486 3732
rect 48682 3720 48688 3732
rect 34992 3692 48688 3720
rect 30374 3612 30380 3664
rect 30432 3652 30438 3664
rect 34701 3655 34759 3661
rect 34701 3652 34713 3655
rect 30432 3624 34713 3652
rect 30432 3612 30438 3624
rect 34701 3621 34713 3624
rect 34747 3621 34759 3655
rect 34701 3615 34759 3621
rect 28074 3544 28080 3596
rect 28132 3584 28138 3596
rect 34992 3584 35020 3692
rect 48682 3680 48688 3692
rect 48740 3680 48746 3732
rect 35066 3612 35072 3664
rect 35124 3612 35130 3664
rect 41601 3655 41659 3661
rect 41601 3621 41613 3655
rect 41647 3652 41659 3655
rect 41782 3652 41788 3664
rect 41647 3624 41788 3652
rect 41647 3621 41659 3624
rect 41601 3615 41659 3621
rect 41782 3612 41788 3624
rect 41840 3612 41846 3664
rect 28132 3556 35020 3584
rect 35084 3584 35112 3612
rect 36449 3587 36507 3593
rect 36449 3584 36461 3587
rect 35084 3556 36461 3584
rect 28132 3544 28138 3556
rect 36449 3553 36461 3556
rect 36495 3553 36507 3587
rect 36449 3547 36507 3553
rect 39853 3587 39911 3593
rect 39853 3553 39865 3587
rect 39899 3584 39911 3587
rect 40218 3584 40224 3596
rect 39899 3556 40224 3584
rect 39899 3553 39911 3556
rect 39853 3547 39911 3553
rect 40218 3544 40224 3556
rect 40276 3544 40282 3596
rect 35158 3408 35164 3460
rect 35216 3408 35222 3460
rect 36173 3451 36231 3457
rect 36173 3417 36185 3451
rect 36219 3417 36231 3451
rect 40126 3448 40132 3460
rect 40087 3420 40132 3448
rect 36173 3411 36231 3417
rect 25424 3352 27752 3380
rect 33042 3340 33048 3392
rect 33100 3380 33106 3392
rect 36188 3380 36216 3411
rect 40126 3408 40132 3420
rect 40184 3408 40190 3460
rect 40402 3408 40408 3460
rect 40460 3448 40466 3460
rect 40460 3420 40618 3448
rect 40460 3408 40466 3420
rect 33100 3352 36216 3380
rect 33100 3340 33106 3352
rect 1104 3290 58880 3312
rect 1104 3238 15398 3290
rect 15450 3238 15462 3290
rect 15514 3238 15526 3290
rect 15578 3238 15590 3290
rect 15642 3238 15654 3290
rect 15706 3238 29846 3290
rect 29898 3238 29910 3290
rect 29962 3238 29974 3290
rect 30026 3238 30038 3290
rect 30090 3238 30102 3290
rect 30154 3238 44294 3290
rect 44346 3238 44358 3290
rect 44410 3238 44422 3290
rect 44474 3238 44486 3290
rect 44538 3238 44550 3290
rect 44602 3238 58880 3290
rect 1104 3216 58880 3238
rect 14185 3179 14243 3185
rect 14185 3145 14197 3179
rect 14231 3176 14243 3179
rect 14274 3176 14280 3188
rect 14231 3148 14280 3176
rect 14231 3145 14243 3148
rect 14185 3139 14243 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 29638 3136 29644 3188
rect 29696 3176 29702 3188
rect 37277 3179 37335 3185
rect 37277 3176 37289 3179
rect 29696 3148 37289 3176
rect 29696 3136 29702 3148
rect 37277 3145 37289 3148
rect 37323 3176 37335 3179
rect 44174 3176 44180 3188
rect 37323 3148 44180 3176
rect 37323 3145 37335 3148
rect 37277 3139 37335 3145
rect 44174 3136 44180 3148
rect 44232 3136 44238 3188
rect 38010 3068 38016 3120
rect 38068 3068 38074 3120
rect 38749 3111 38807 3117
rect 38749 3077 38761 3111
rect 38795 3108 38807 3111
rect 41230 3108 41236 3120
rect 38795 3080 41236 3108
rect 38795 3077 38807 3080
rect 38749 3071 38807 3077
rect 41230 3068 41236 3080
rect 41288 3068 41294 3120
rect 19702 3000 19708 3052
rect 19760 3040 19766 3052
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19760 3012 19809 3040
rect 19760 3000 19766 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 27890 3040 27896 3052
rect 27851 3012 27896 3040
rect 19797 3003 19855 3009
rect 27890 3000 27896 3012
rect 27948 3040 27954 3052
rect 28537 3043 28595 3049
rect 28537 3040 28549 3043
rect 27948 3012 28549 3040
rect 27948 3000 27954 3012
rect 28537 3009 28549 3012
rect 28583 3009 28595 3043
rect 28537 3003 28595 3009
rect 32398 3000 32404 3052
rect 32456 3040 32462 3052
rect 33321 3043 33379 3049
rect 33321 3040 33333 3043
rect 32456 3012 33333 3040
rect 32456 3000 32462 3012
rect 33321 3009 33333 3012
rect 33367 3040 33379 3043
rect 34882 3040 34888 3052
rect 33367 3012 34888 3040
rect 33367 3009 33379 3012
rect 33321 3003 33379 3009
rect 34882 3000 34888 3012
rect 34940 3000 34946 3052
rect 48866 3000 48872 3052
rect 48924 3040 48930 3052
rect 57885 3043 57943 3049
rect 57885 3040 57897 3043
rect 48924 3012 57897 3040
rect 48924 3000 48930 3012
rect 57885 3009 57897 3012
rect 57931 3009 57943 3043
rect 57885 3003 57943 3009
rect 29178 2932 29184 2984
rect 29236 2972 29242 2984
rect 39025 2975 39083 2981
rect 29236 2944 37228 2972
rect 29236 2932 29242 2944
rect 28077 2907 28135 2913
rect 28077 2873 28089 2907
rect 28123 2904 28135 2907
rect 29546 2904 29552 2916
rect 28123 2876 29552 2904
rect 28123 2873 28135 2876
rect 28077 2867 28135 2873
rect 29546 2864 29552 2876
rect 29604 2864 29610 2916
rect 19613 2839 19671 2845
rect 19613 2805 19625 2839
rect 19659 2836 19671 2839
rect 19702 2836 19708 2848
rect 19659 2808 19708 2836
rect 19659 2805 19671 2808
rect 19613 2799 19671 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 33505 2839 33563 2845
rect 33505 2805 33517 2839
rect 33551 2836 33563 2839
rect 33778 2836 33784 2848
rect 33551 2808 33784 2836
rect 33551 2805 33563 2808
rect 33505 2799 33563 2805
rect 33778 2796 33784 2808
rect 33836 2796 33842 2848
rect 37200 2836 37228 2944
rect 39025 2941 39037 2975
rect 39071 2972 39083 2975
rect 39485 2975 39543 2981
rect 39485 2972 39497 2975
rect 39071 2944 39497 2972
rect 39071 2941 39083 2944
rect 39025 2935 39083 2941
rect 39485 2941 39497 2944
rect 39531 2972 39543 2975
rect 39531 2944 41414 2972
rect 39531 2941 39543 2944
rect 39485 2935 39543 2941
rect 39040 2836 39068 2935
rect 41386 2904 41414 2944
rect 53098 2904 53104 2916
rect 41386 2876 53104 2904
rect 53098 2864 53104 2876
rect 53156 2864 53162 2916
rect 37200 2808 39068 2836
rect 52822 2796 52828 2848
rect 52880 2836 52886 2848
rect 52917 2839 52975 2845
rect 52917 2836 52929 2839
rect 52880 2808 52929 2836
rect 52880 2796 52886 2808
rect 52917 2805 52929 2808
rect 52963 2805 52975 2839
rect 58066 2836 58072 2848
rect 58027 2808 58072 2836
rect 52917 2799 52975 2805
rect 58066 2796 58072 2808
rect 58124 2796 58130 2848
rect 1104 2746 58880 2768
rect 1104 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 8302 2746
rect 8354 2694 8366 2746
rect 8418 2694 8430 2746
rect 8482 2694 22622 2746
rect 22674 2694 22686 2746
rect 22738 2694 22750 2746
rect 22802 2694 22814 2746
rect 22866 2694 22878 2746
rect 22930 2694 37070 2746
rect 37122 2694 37134 2746
rect 37186 2694 37198 2746
rect 37250 2694 37262 2746
rect 37314 2694 37326 2746
rect 37378 2694 51518 2746
rect 51570 2694 51582 2746
rect 51634 2694 51646 2746
rect 51698 2694 51710 2746
rect 51762 2694 51774 2746
rect 51826 2694 58880 2746
rect 1104 2672 58880 2694
rect 37826 2592 37832 2644
rect 37884 2632 37890 2644
rect 38197 2635 38255 2641
rect 38197 2632 38209 2635
rect 37884 2604 38209 2632
rect 37884 2592 37890 2604
rect 38197 2601 38209 2604
rect 38243 2601 38255 2635
rect 38197 2595 38255 2601
rect 10045 2567 10103 2573
rect 10045 2533 10057 2567
rect 10091 2564 10103 2567
rect 13814 2564 13820 2576
rect 10091 2536 13820 2564
rect 10091 2533 10103 2536
rect 10045 2527 10103 2533
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4522 2428 4528 2440
rect 4203 2400 4528 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 4522 2388 4528 2400
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 14274 2428 14280 2440
rect 14235 2400 14280 2428
rect 4617 2391 4675 2397
rect 14274 2388 14280 2400
rect 14332 2388 14338 2440
rect 19702 2428 19708 2440
rect 19663 2400 19708 2428
rect 19702 2388 19708 2400
rect 19760 2388 19766 2440
rect 24673 2431 24731 2437
rect 24673 2397 24685 2431
rect 24719 2397 24731 2431
rect 29546 2428 29552 2440
rect 29507 2400 29552 2428
rect 24673 2391 24731 2397
rect 9309 2363 9367 2369
rect 9309 2329 9321 2363
rect 9355 2360 9367 2363
rect 9674 2360 9680 2372
rect 9355 2332 9680 2360
rect 9355 2329 9367 2332
rect 9309 2323 9367 2329
rect 9674 2320 9680 2332
rect 9732 2360 9738 2372
rect 9861 2363 9919 2369
rect 9861 2360 9873 2363
rect 9732 2332 9873 2360
rect 9732 2320 9738 2332
rect 9861 2329 9873 2332
rect 9907 2329 9919 2363
rect 16298 2360 16304 2372
rect 9861 2323 9919 2329
rect 11256 2332 16304 2360
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1489 2295 1547 2301
rect 1489 2292 1501 2295
rect 72 2264 1501 2292
rect 72 2252 78 2264
rect 1489 2261 1501 2264
rect 1535 2261 1547 2295
rect 1489 2255 1547 2261
rect 4801 2295 4859 2301
rect 4801 2261 4813 2295
rect 4847 2292 4859 2295
rect 11256 2292 11284 2332
rect 16298 2320 16304 2332
rect 16356 2320 16362 2372
rect 24688 2360 24716 2391
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 33778 2428 33784 2440
rect 33739 2400 33784 2428
rect 33778 2388 33784 2400
rect 33836 2388 33842 2440
rect 38212 2428 38240 2595
rect 41230 2592 41236 2644
rect 41288 2632 41294 2644
rect 43257 2635 43315 2641
rect 43257 2632 43269 2635
rect 41288 2604 43269 2632
rect 41288 2592 41294 2604
rect 43257 2601 43269 2604
rect 43303 2601 43315 2635
rect 43257 2595 43315 2601
rect 53098 2564 53104 2576
rect 53059 2536 53104 2564
rect 53098 2524 53104 2536
rect 53156 2524 53162 2576
rect 38749 2431 38807 2437
rect 38749 2428 38761 2431
rect 38212 2400 38761 2428
rect 38749 2397 38761 2400
rect 38795 2397 38807 2431
rect 38749 2391 38807 2397
rect 43162 2388 43168 2440
rect 43220 2428 43226 2440
rect 43441 2431 43499 2437
rect 43441 2428 43453 2431
rect 43220 2400 43453 2428
rect 43220 2388 43226 2400
rect 43441 2397 43453 2400
rect 43487 2428 43499 2431
rect 43901 2431 43959 2437
rect 43901 2428 43913 2431
rect 43487 2400 43913 2428
rect 43487 2397 43499 2400
rect 43441 2391 43499 2397
rect 43901 2397 43913 2400
rect 43947 2397 43959 2431
rect 48406 2428 48412 2440
rect 48367 2400 48412 2428
rect 43901 2391 43959 2397
rect 48406 2388 48412 2400
rect 48464 2388 48470 2440
rect 57882 2428 57888 2440
rect 57843 2400 57888 2428
rect 57882 2388 57888 2400
rect 57940 2388 57946 2440
rect 25225 2363 25283 2369
rect 25225 2360 25237 2363
rect 24688 2332 25237 2360
rect 25225 2329 25237 2332
rect 25271 2360 25283 2363
rect 41414 2360 41420 2372
rect 25271 2332 41420 2360
rect 25271 2329 25283 2332
rect 25225 2323 25283 2329
rect 41414 2320 41420 2332
rect 41472 2320 41478 2372
rect 52822 2320 52828 2372
rect 52880 2360 52886 2372
rect 53285 2363 53343 2369
rect 53285 2360 53297 2363
rect 52880 2332 53297 2360
rect 52880 2320 52886 2332
rect 53285 2329 53297 2332
rect 53331 2329 53343 2363
rect 53285 2323 53343 2329
rect 4847 2264 11284 2292
rect 4847 2261 4859 2264
rect 4801 2255 4859 2261
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 14240 2264 14473 2292
rect 14240 2252 14246 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19521 2295 19579 2301
rect 19521 2292 19533 2295
rect 19392 2264 19533 2292
rect 19392 2252 19398 2264
rect 19521 2261 19533 2264
rect 19567 2261 19579 2295
rect 19521 2255 19579 2261
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24489 2295 24547 2301
rect 24489 2292 24501 2295
rect 23900 2264 24501 2292
rect 23900 2252 23906 2264
rect 24489 2261 24501 2264
rect 24535 2261 24547 2295
rect 24489 2255 24547 2261
rect 28994 2252 29000 2304
rect 29052 2292 29058 2304
rect 29733 2295 29791 2301
rect 29733 2292 29745 2295
rect 29052 2264 29745 2292
rect 29052 2252 29058 2264
rect 29733 2261 29745 2264
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33597 2295 33655 2301
rect 33597 2292 33609 2295
rect 33560 2264 33609 2292
rect 33560 2252 33566 2264
rect 33597 2261 33609 2264
rect 33643 2261 33655 2295
rect 33597 2255 33655 2261
rect 38654 2252 38660 2304
rect 38712 2292 38718 2304
rect 38933 2295 38991 2301
rect 38933 2292 38945 2295
rect 38712 2264 38945 2292
rect 38712 2252 38718 2264
rect 38933 2261 38945 2264
rect 38979 2261 38991 2295
rect 38933 2255 38991 2261
rect 48314 2252 48320 2304
rect 48372 2292 48378 2304
rect 48593 2295 48651 2301
rect 48593 2292 48605 2295
rect 48372 2264 48605 2292
rect 48372 2252 48378 2264
rect 48593 2261 48605 2264
rect 48639 2261 48651 2295
rect 48593 2255 48651 2261
rect 57974 2252 57980 2304
rect 58032 2292 58038 2304
rect 58069 2295 58127 2301
rect 58069 2292 58081 2295
rect 58032 2264 58081 2292
rect 58032 2252 58038 2264
rect 58069 2261 58081 2264
rect 58115 2261 58127 2295
rect 58069 2255 58127 2261
rect 1104 2202 58880 2224
rect 1104 2150 15398 2202
rect 15450 2150 15462 2202
rect 15514 2150 15526 2202
rect 15578 2150 15590 2202
rect 15642 2150 15654 2202
rect 15706 2150 29846 2202
rect 29898 2150 29910 2202
rect 29962 2150 29974 2202
rect 30026 2150 30038 2202
rect 30090 2150 30102 2202
rect 30154 2150 44294 2202
rect 44346 2150 44358 2202
rect 44410 2150 44422 2202
rect 44474 2150 44486 2202
rect 44538 2150 44550 2202
rect 44602 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 15398 33702 15450 33754
rect 15462 33702 15514 33754
rect 15526 33702 15578 33754
rect 15590 33702 15642 33754
rect 15654 33702 15706 33754
rect 29846 33702 29898 33754
rect 29910 33702 29962 33754
rect 29974 33702 30026 33754
rect 30038 33702 30090 33754
rect 30102 33702 30154 33754
rect 44294 33702 44346 33754
rect 44358 33702 44410 33754
rect 44422 33702 44474 33754
rect 44486 33702 44538 33754
rect 44550 33702 44602 33754
rect 1492 33643 1544 33652
rect 1492 33609 1501 33643
rect 1501 33609 1535 33643
rect 1535 33609 1544 33643
rect 1492 33600 1544 33609
rect 4804 33643 4856 33652
rect 4804 33609 4813 33643
rect 4813 33609 4847 33643
rect 4847 33609 4856 33643
rect 4804 33600 4856 33609
rect 9036 33600 9088 33652
rect 14372 33643 14424 33652
rect 14372 33609 14381 33643
rect 14381 33609 14415 33643
rect 14415 33609 14424 33643
rect 14372 33600 14424 33609
rect 18696 33600 18748 33652
rect 33784 33643 33836 33652
rect 33784 33609 33793 33643
rect 33793 33609 33827 33643
rect 33827 33609 33836 33643
rect 33784 33600 33836 33609
rect 38660 33600 38712 33652
rect 43260 33643 43312 33652
rect 43260 33609 43269 33643
rect 43269 33609 43303 33643
rect 43303 33609 43312 33643
rect 43260 33600 43312 33609
rect 48596 33643 48648 33652
rect 48596 33609 48605 33643
rect 48605 33609 48639 33643
rect 48639 33609 48648 33643
rect 48596 33600 48648 33609
rect 53104 33643 53156 33652
rect 53104 33609 53113 33643
rect 53113 33609 53147 33643
rect 53147 33609 53156 33643
rect 53104 33600 53156 33609
rect 28540 33575 28592 33584
rect 28540 33541 28549 33575
rect 28549 33541 28583 33575
rect 28583 33541 28592 33575
rect 28540 33532 28592 33541
rect 1676 33507 1728 33516
rect 1676 33473 1685 33507
rect 1685 33473 1719 33507
rect 1719 33473 1728 33507
rect 1676 33464 1728 33473
rect 4620 33507 4672 33516
rect 4620 33473 4629 33507
rect 4629 33473 4663 33507
rect 4663 33473 4672 33507
rect 4620 33464 4672 33473
rect 9404 33507 9456 33516
rect 9404 33473 9413 33507
rect 9413 33473 9447 33507
rect 9447 33473 9456 33507
rect 9404 33464 9456 33473
rect 17224 33464 17276 33516
rect 19432 33507 19484 33516
rect 19432 33473 19441 33507
rect 19441 33473 19475 33507
rect 19475 33473 19484 33507
rect 19432 33464 19484 33473
rect 23848 33464 23900 33516
rect 6828 33260 6880 33312
rect 8024 33260 8076 33312
rect 24400 33303 24452 33312
rect 24400 33269 24409 33303
rect 24409 33269 24443 33303
rect 24443 33269 24452 33303
rect 24400 33260 24452 33269
rect 27344 33260 27396 33312
rect 33600 33507 33652 33516
rect 33600 33473 33609 33507
rect 33609 33473 33643 33507
rect 33643 33473 33652 33507
rect 33600 33464 33652 33473
rect 38936 33507 38988 33516
rect 38936 33473 38945 33507
rect 38945 33473 38979 33507
rect 38979 33473 38988 33507
rect 38936 33464 38988 33473
rect 43904 33464 43956 33516
rect 48412 33507 48464 33516
rect 48412 33473 48421 33507
rect 48421 33473 48455 33507
rect 48455 33473 48464 33507
rect 48412 33464 48464 33473
rect 52644 33464 52696 33516
rect 57796 33464 57848 33516
rect 56600 33396 56652 33448
rect 36268 33328 36320 33380
rect 58072 33371 58124 33380
rect 58072 33337 58081 33371
rect 58081 33337 58115 33371
rect 58115 33337 58124 33371
rect 58072 33328 58124 33337
rect 35900 33303 35952 33312
rect 35900 33269 35909 33303
rect 35909 33269 35943 33303
rect 35943 33269 35952 33303
rect 35900 33260 35952 33269
rect 37740 33260 37792 33312
rect 57520 33260 57572 33312
rect 8174 33158 8226 33210
rect 8238 33158 8290 33210
rect 8302 33158 8354 33210
rect 8366 33158 8418 33210
rect 8430 33158 8482 33210
rect 22622 33158 22674 33210
rect 22686 33158 22738 33210
rect 22750 33158 22802 33210
rect 22814 33158 22866 33210
rect 22878 33158 22930 33210
rect 37070 33158 37122 33210
rect 37134 33158 37186 33210
rect 37198 33158 37250 33210
rect 37262 33158 37314 33210
rect 37326 33158 37378 33210
rect 51518 33158 51570 33210
rect 51582 33158 51634 33210
rect 51646 33158 51698 33210
rect 51710 33158 51762 33210
rect 51774 33158 51826 33210
rect 4620 33056 4672 33108
rect 19432 33099 19484 33108
rect 19432 33065 19441 33099
rect 19441 33065 19475 33099
rect 19475 33065 19484 33099
rect 19432 33056 19484 33065
rect 33600 33056 33652 33108
rect 38936 33056 38988 33108
rect 57796 33056 57848 33108
rect 4436 32852 4488 32904
rect 5172 32895 5224 32904
rect 5172 32861 5181 32895
rect 5181 32861 5215 32895
rect 5215 32861 5224 32895
rect 5172 32852 5224 32861
rect 5448 32895 5500 32904
rect 5448 32861 5457 32895
rect 5457 32861 5491 32895
rect 5491 32861 5500 32895
rect 5448 32852 5500 32861
rect 6552 32852 6604 32904
rect 18696 32895 18748 32904
rect 18696 32861 18705 32895
rect 18705 32861 18739 32895
rect 18739 32861 18748 32895
rect 18696 32852 18748 32861
rect 6920 32784 6972 32836
rect 6368 32759 6420 32768
rect 6368 32725 6377 32759
rect 6377 32725 6411 32759
rect 6411 32725 6420 32759
rect 6368 32716 6420 32725
rect 7012 32716 7064 32768
rect 9404 32716 9456 32768
rect 35808 32852 35860 32904
rect 36452 32852 36504 32904
rect 37740 32895 37792 32904
rect 37740 32861 37749 32895
rect 37749 32861 37783 32895
rect 37783 32861 37792 32895
rect 37740 32852 37792 32861
rect 24308 32716 24360 32768
rect 32956 32759 33008 32768
rect 32956 32725 32965 32759
rect 32965 32725 32999 32759
rect 32999 32725 33008 32759
rect 32956 32716 33008 32725
rect 35716 32716 35768 32768
rect 37556 32784 37608 32836
rect 48412 32716 48464 32768
rect 52644 32716 52696 32768
rect 15398 32614 15450 32666
rect 15462 32614 15514 32666
rect 15526 32614 15578 32666
rect 15590 32614 15642 32666
rect 15654 32614 15706 32666
rect 29846 32614 29898 32666
rect 29910 32614 29962 32666
rect 29974 32614 30026 32666
rect 30038 32614 30090 32666
rect 30102 32614 30154 32666
rect 44294 32614 44346 32666
rect 44358 32614 44410 32666
rect 44422 32614 44474 32666
rect 44486 32614 44538 32666
rect 44550 32614 44602 32666
rect 6552 32555 6604 32564
rect 6552 32521 6561 32555
rect 6561 32521 6595 32555
rect 6595 32521 6604 32555
rect 6552 32512 6604 32521
rect 37740 32512 37792 32564
rect 38568 32512 38620 32564
rect 5448 32444 5500 32496
rect 2780 32419 2832 32428
rect 2780 32385 2789 32419
rect 2789 32385 2823 32419
rect 2823 32385 2832 32419
rect 2780 32376 2832 32385
rect 7012 32444 7064 32496
rect 7932 32444 7984 32496
rect 36268 32444 36320 32496
rect 1768 32351 1820 32360
rect 1768 32317 1777 32351
rect 1777 32317 1811 32351
rect 1811 32317 1820 32351
rect 1768 32308 1820 32317
rect 6920 32308 6972 32360
rect 9036 32351 9088 32360
rect 3056 32172 3108 32224
rect 4436 32172 4488 32224
rect 9036 32317 9045 32351
rect 9045 32317 9079 32351
rect 9079 32317 9088 32351
rect 9036 32308 9088 32317
rect 24400 32172 24452 32224
rect 35716 32215 35768 32224
rect 35716 32181 35725 32215
rect 35725 32181 35759 32215
rect 35759 32181 35768 32215
rect 35716 32172 35768 32181
rect 35808 32172 35860 32224
rect 37464 32215 37516 32224
rect 37464 32181 37473 32215
rect 37473 32181 37507 32215
rect 37507 32181 37516 32215
rect 37464 32172 37516 32181
rect 37924 32172 37976 32224
rect 38476 32172 38528 32224
rect 8174 32070 8226 32122
rect 8238 32070 8290 32122
rect 8302 32070 8354 32122
rect 8366 32070 8418 32122
rect 8430 32070 8482 32122
rect 22622 32070 22674 32122
rect 22686 32070 22738 32122
rect 22750 32070 22802 32122
rect 22814 32070 22866 32122
rect 22878 32070 22930 32122
rect 37070 32070 37122 32122
rect 37134 32070 37186 32122
rect 37198 32070 37250 32122
rect 37262 32070 37314 32122
rect 37326 32070 37378 32122
rect 51518 32070 51570 32122
rect 51582 32070 51634 32122
rect 51646 32070 51698 32122
rect 51710 32070 51762 32122
rect 51774 32070 51826 32122
rect 37556 31968 37608 32020
rect 38568 31968 38620 32020
rect 8024 31875 8076 31884
rect 8024 31841 8033 31875
rect 8033 31841 8067 31875
rect 8067 31841 8076 31875
rect 8024 31832 8076 31841
rect 1768 31764 1820 31816
rect 5172 31807 5224 31816
rect 5172 31773 5181 31807
rect 5181 31773 5215 31807
rect 5215 31773 5224 31807
rect 5172 31764 5224 31773
rect 5448 31807 5500 31816
rect 5448 31773 5457 31807
rect 5457 31773 5491 31807
rect 5491 31773 5500 31807
rect 5448 31764 5500 31773
rect 6184 31807 6236 31816
rect 6184 31773 6193 31807
rect 6193 31773 6227 31807
rect 6227 31773 6236 31807
rect 6184 31764 6236 31773
rect 6552 31764 6604 31816
rect 4620 31671 4672 31680
rect 4620 31637 4629 31671
rect 4629 31637 4663 31671
rect 4663 31637 4672 31671
rect 4620 31628 4672 31637
rect 6368 31671 6420 31680
rect 6368 31637 6377 31671
rect 6377 31637 6411 31671
rect 6411 31637 6420 31671
rect 6368 31628 6420 31637
rect 7656 31628 7708 31680
rect 35164 31628 35216 31680
rect 35808 31764 35860 31816
rect 35716 31696 35768 31748
rect 37464 31764 37516 31816
rect 37924 31807 37976 31816
rect 37924 31773 37933 31807
rect 37933 31773 37967 31807
rect 37967 31773 37976 31807
rect 37924 31764 37976 31773
rect 38476 31764 38528 31816
rect 15398 31526 15450 31578
rect 15462 31526 15514 31578
rect 15526 31526 15578 31578
rect 15590 31526 15642 31578
rect 15654 31526 15706 31578
rect 29846 31526 29898 31578
rect 29910 31526 29962 31578
rect 29974 31526 30026 31578
rect 30038 31526 30090 31578
rect 30102 31526 30154 31578
rect 44294 31526 44346 31578
rect 44358 31526 44410 31578
rect 44422 31526 44474 31578
rect 44486 31526 44538 31578
rect 44550 31526 44602 31578
rect 37556 31424 37608 31476
rect 38476 31424 38528 31476
rect 3056 31356 3108 31408
rect 5816 31399 5868 31408
rect 5816 31365 5825 31399
rect 5825 31365 5859 31399
rect 5859 31365 5868 31399
rect 6368 31399 6420 31408
rect 5816 31356 5868 31365
rect 6368 31365 6377 31399
rect 6377 31365 6411 31399
rect 6411 31365 6420 31399
rect 6368 31356 6420 31365
rect 5448 31288 5500 31340
rect 6184 31288 6236 31340
rect 7656 31288 7708 31340
rect 35716 31288 35768 31340
rect 37464 31331 37516 31340
rect 37464 31297 37473 31331
rect 37473 31297 37507 31331
rect 37507 31297 37516 31331
rect 37464 31288 37516 31297
rect 38568 31288 38620 31340
rect 45836 31331 45888 31340
rect 45836 31297 45845 31331
rect 45845 31297 45879 31331
rect 45879 31297 45888 31331
rect 45836 31288 45888 31297
rect 8024 31220 8076 31272
rect 35164 31220 35216 31272
rect 4620 31084 4672 31136
rect 7656 31084 7708 31136
rect 56600 31084 56652 31136
rect 8174 30982 8226 31034
rect 8238 30982 8290 31034
rect 8302 30982 8354 31034
rect 8366 30982 8418 31034
rect 8430 30982 8482 31034
rect 22622 30982 22674 31034
rect 22686 30982 22738 31034
rect 22750 30982 22802 31034
rect 22814 30982 22866 31034
rect 22878 30982 22930 31034
rect 37070 30982 37122 31034
rect 37134 30982 37186 31034
rect 37198 30982 37250 31034
rect 37262 30982 37314 31034
rect 37326 30982 37378 31034
rect 51518 30982 51570 31034
rect 51582 30982 51634 31034
rect 51646 30982 51698 31034
rect 51710 30982 51762 31034
rect 51774 30982 51826 31034
rect 1676 30880 1728 30932
rect 5816 30880 5868 30932
rect 6828 30923 6880 30932
rect 6828 30889 6837 30923
rect 6837 30889 6871 30923
rect 6871 30889 6880 30923
rect 6828 30880 6880 30889
rect 37556 30880 37608 30932
rect 38568 30880 38620 30932
rect 2872 30676 2924 30728
rect 3056 30719 3108 30728
rect 3056 30685 3065 30719
rect 3065 30685 3099 30719
rect 3099 30685 3108 30719
rect 3056 30676 3108 30685
rect 4620 30676 4672 30728
rect 5448 30719 5500 30728
rect 5448 30685 5457 30719
rect 5457 30685 5491 30719
rect 5491 30685 5500 30719
rect 5448 30676 5500 30685
rect 6184 30719 6236 30728
rect 6184 30685 6193 30719
rect 6193 30685 6227 30719
rect 6227 30685 6236 30719
rect 6184 30676 6236 30685
rect 6552 30676 6604 30728
rect 8024 30719 8076 30728
rect 1492 30583 1544 30592
rect 1492 30549 1501 30583
rect 1501 30549 1535 30583
rect 1535 30549 1544 30583
rect 1492 30540 1544 30549
rect 4620 30583 4672 30592
rect 4620 30549 4629 30583
rect 4629 30549 4663 30583
rect 4663 30549 4672 30583
rect 4620 30540 4672 30549
rect 7656 30540 7708 30592
rect 8024 30685 8033 30719
rect 8033 30685 8067 30719
rect 8067 30685 8076 30719
rect 8024 30676 8076 30685
rect 35808 30676 35860 30728
rect 37464 30676 37516 30728
rect 37924 30719 37976 30728
rect 37924 30685 37933 30719
rect 37933 30685 37967 30719
rect 37967 30685 37976 30719
rect 37924 30676 37976 30685
rect 38476 30676 38528 30728
rect 35164 30540 35216 30592
rect 35348 30540 35400 30592
rect 37372 30608 37424 30660
rect 15398 30438 15450 30490
rect 15462 30438 15514 30490
rect 15526 30438 15578 30490
rect 15590 30438 15642 30490
rect 15654 30438 15706 30490
rect 29846 30438 29898 30490
rect 29910 30438 29962 30490
rect 29974 30438 30026 30490
rect 30038 30438 30090 30490
rect 30102 30438 30154 30490
rect 44294 30438 44346 30490
rect 44358 30438 44410 30490
rect 44422 30438 44474 30490
rect 44486 30438 44538 30490
rect 44550 30438 44602 30490
rect 5816 30379 5868 30388
rect 5816 30345 5825 30379
rect 5825 30345 5859 30379
rect 5859 30345 5868 30379
rect 5816 30336 5868 30345
rect 6184 30336 6236 30388
rect 37372 30336 37424 30388
rect 38476 30336 38528 30388
rect 5448 30200 5500 30252
rect 7012 30268 7064 30320
rect 6552 30200 6604 30252
rect 6828 30200 6880 30252
rect 7840 30200 7892 30252
rect 14372 30200 14424 30252
rect 19524 30243 19576 30252
rect 19524 30209 19533 30243
rect 19533 30209 19567 30243
rect 19567 30209 19576 30243
rect 19524 30200 19576 30209
rect 4620 30175 4672 30184
rect 4620 30141 4629 30175
rect 4629 30141 4663 30175
rect 4663 30141 4672 30175
rect 4620 30132 4672 30141
rect 14556 30132 14608 30184
rect 4160 30039 4212 30048
rect 4160 30005 4169 30039
rect 4169 30005 4203 30039
rect 4203 30005 4212 30039
rect 4160 29996 4212 30005
rect 7656 30039 7708 30048
rect 7656 30005 7665 30039
rect 7665 30005 7699 30039
rect 7699 30005 7708 30039
rect 7656 29996 7708 30005
rect 8024 29996 8076 30048
rect 15200 30039 15252 30048
rect 15200 30005 15209 30039
rect 15209 30005 15243 30039
rect 15243 30005 15252 30039
rect 15200 29996 15252 30005
rect 20720 29996 20772 30048
rect 35808 29996 35860 30048
rect 8174 29894 8226 29946
rect 8238 29894 8290 29946
rect 8302 29894 8354 29946
rect 8366 29894 8418 29946
rect 8430 29894 8482 29946
rect 22622 29894 22674 29946
rect 22686 29894 22738 29946
rect 22750 29894 22802 29946
rect 22814 29894 22866 29946
rect 22878 29894 22930 29946
rect 37070 29894 37122 29946
rect 37134 29894 37186 29946
rect 37198 29894 37250 29946
rect 37262 29894 37314 29946
rect 37326 29894 37378 29946
rect 51518 29894 51570 29946
rect 51582 29894 51634 29946
rect 51646 29894 51698 29946
rect 51710 29894 51762 29946
rect 51774 29894 51826 29946
rect 15200 29792 15252 29844
rect 2504 29656 2556 29708
rect 6920 29724 6972 29776
rect 4068 29563 4120 29572
rect 4068 29529 4077 29563
rect 4077 29529 4111 29563
rect 4111 29529 4120 29563
rect 4068 29520 4120 29529
rect 3240 29452 3292 29504
rect 14556 29699 14608 29708
rect 14556 29665 14565 29699
rect 14565 29665 14599 29699
rect 14599 29665 14608 29699
rect 14556 29656 14608 29665
rect 19524 29656 19576 29708
rect 20720 29699 20772 29708
rect 20720 29665 20729 29699
rect 20729 29665 20763 29699
rect 20763 29665 20772 29699
rect 20720 29656 20772 29665
rect 37556 29792 37608 29844
rect 27528 29656 27580 29708
rect 6000 29631 6052 29640
rect 6000 29597 6009 29631
rect 6009 29597 6043 29631
rect 6043 29597 6052 29631
rect 6000 29588 6052 29597
rect 14372 29588 14424 29640
rect 7012 29520 7064 29572
rect 16488 29563 16540 29572
rect 16488 29529 16497 29563
rect 16497 29529 16531 29563
rect 16531 29529 16540 29563
rect 16488 29520 16540 29529
rect 18604 29563 18656 29572
rect 5356 29452 5408 29504
rect 6276 29452 6328 29504
rect 8024 29452 8076 29504
rect 9588 29452 9640 29504
rect 15752 29495 15804 29504
rect 15752 29461 15761 29495
rect 15761 29461 15795 29495
rect 15795 29461 15804 29495
rect 18604 29529 18613 29563
rect 18613 29529 18647 29563
rect 18647 29529 18656 29563
rect 18604 29520 18656 29529
rect 20628 29520 20680 29572
rect 24124 29588 24176 29640
rect 35164 29588 35216 29640
rect 35808 29588 35860 29640
rect 27160 29563 27212 29572
rect 27160 29529 27169 29563
rect 27169 29529 27203 29563
rect 27203 29529 27212 29563
rect 27160 29520 27212 29529
rect 37924 29588 37976 29640
rect 19248 29495 19300 29504
rect 15752 29452 15804 29461
rect 19248 29461 19257 29495
rect 19257 29461 19291 29495
rect 19291 29461 19300 29495
rect 19248 29452 19300 29461
rect 26424 29495 26476 29504
rect 26424 29461 26433 29495
rect 26433 29461 26467 29495
rect 26467 29461 26476 29495
rect 26424 29452 26476 29461
rect 30196 29452 30248 29504
rect 35348 29452 35400 29504
rect 15398 29350 15450 29402
rect 15462 29350 15514 29402
rect 15526 29350 15578 29402
rect 15590 29350 15642 29402
rect 15654 29350 15706 29402
rect 29846 29350 29898 29402
rect 29910 29350 29962 29402
rect 29974 29350 30026 29402
rect 30038 29350 30090 29402
rect 30102 29350 30154 29402
rect 44294 29350 44346 29402
rect 44358 29350 44410 29402
rect 44422 29350 44474 29402
rect 44486 29350 44538 29402
rect 44550 29350 44602 29402
rect 4068 29248 4120 29300
rect 7012 29248 7064 29300
rect 16488 29248 16540 29300
rect 24124 29291 24176 29300
rect 24124 29257 24133 29291
rect 24133 29257 24167 29291
rect 24167 29257 24176 29291
rect 24124 29248 24176 29257
rect 2780 29180 2832 29232
rect 3240 29180 3292 29232
rect 4160 29180 4212 29232
rect 6736 29180 6788 29232
rect 2504 29155 2556 29164
rect 2504 29121 2513 29155
rect 2513 29121 2547 29155
rect 2547 29121 2556 29155
rect 2504 29112 2556 29121
rect 7012 29044 7064 29096
rect 8024 29044 8076 29096
rect 19248 29112 19300 29164
rect 26424 29180 26476 29232
rect 19524 29044 19576 29096
rect 21732 29044 21784 29096
rect 26792 29112 26844 29164
rect 36268 29155 36320 29164
rect 36268 29121 36277 29155
rect 36277 29121 36311 29155
rect 36311 29121 36320 29155
rect 36268 29112 36320 29121
rect 27528 29087 27580 29096
rect 27528 29053 27537 29087
rect 27537 29053 27571 29087
rect 27571 29053 27580 29087
rect 27528 29044 27580 29053
rect 28908 29044 28960 29096
rect 5356 29019 5408 29028
rect 5356 28985 5365 29019
rect 5365 28985 5399 29019
rect 5399 28985 5408 29019
rect 5356 28976 5408 28985
rect 6184 28976 6236 29028
rect 8760 29019 8812 29028
rect 8760 28985 8769 29019
rect 8769 28985 8803 29019
rect 8803 28985 8812 29019
rect 8760 28976 8812 28985
rect 36084 29019 36136 29028
rect 36084 28985 36093 29019
rect 36093 28985 36127 29019
rect 36127 28985 36136 29019
rect 36084 28976 36136 28985
rect 2320 28908 2372 28960
rect 4988 28908 5040 28960
rect 6368 28908 6420 28960
rect 18052 28908 18104 28960
rect 27436 28908 27488 28960
rect 34796 28951 34848 28960
rect 34796 28917 34805 28951
rect 34805 28917 34839 28951
rect 34839 28917 34848 28951
rect 34796 28908 34848 28917
rect 8174 28806 8226 28858
rect 8238 28806 8290 28858
rect 8302 28806 8354 28858
rect 8366 28806 8418 28858
rect 8430 28806 8482 28858
rect 22622 28806 22674 28858
rect 22686 28806 22738 28858
rect 22750 28806 22802 28858
rect 22814 28806 22866 28858
rect 22878 28806 22930 28858
rect 37070 28806 37122 28858
rect 37134 28806 37186 28858
rect 37198 28806 37250 28858
rect 37262 28806 37314 28858
rect 37326 28806 37378 28858
rect 51518 28806 51570 28858
rect 51582 28806 51634 28858
rect 51646 28806 51698 28858
rect 51710 28806 51762 28858
rect 51774 28806 51826 28858
rect 6000 28704 6052 28756
rect 7840 28704 7892 28756
rect 18604 28747 18656 28756
rect 18604 28713 18613 28747
rect 18613 28713 18647 28747
rect 18647 28713 18656 28747
rect 18604 28704 18656 28713
rect 27160 28704 27212 28756
rect 27436 28747 27488 28756
rect 27436 28713 27445 28747
rect 27445 28713 27479 28747
rect 27479 28713 27488 28747
rect 27436 28704 27488 28713
rect 37556 28704 37608 28756
rect 4988 28636 5040 28688
rect 9680 28568 9732 28620
rect 14556 28568 14608 28620
rect 5356 28500 5408 28552
rect 6184 28543 6236 28552
rect 6184 28509 6193 28543
rect 6193 28509 6227 28543
rect 6227 28509 6236 28543
rect 6184 28500 6236 28509
rect 6276 28500 6328 28552
rect 6736 28500 6788 28552
rect 7012 28543 7064 28552
rect 7012 28509 7021 28543
rect 7021 28509 7055 28543
rect 7055 28509 7064 28543
rect 7012 28500 7064 28509
rect 7932 28543 7984 28552
rect 4344 28432 4396 28484
rect 7932 28509 7941 28543
rect 7941 28509 7975 28543
rect 7975 28509 7984 28543
rect 7932 28500 7984 28509
rect 14372 28543 14424 28552
rect 14372 28509 14381 28543
rect 14381 28509 14415 28543
rect 14415 28509 14424 28543
rect 14372 28500 14424 28509
rect 17776 28500 17828 28552
rect 26792 28543 26844 28552
rect 26792 28509 26801 28543
rect 26801 28509 26835 28543
rect 26835 28509 26844 28543
rect 26792 28500 26844 28509
rect 27528 28543 27580 28552
rect 27528 28509 27537 28543
rect 27537 28509 27571 28543
rect 27571 28509 27580 28543
rect 27528 28500 27580 28509
rect 35348 28543 35400 28552
rect 7656 28432 7708 28484
rect 6460 28364 6512 28416
rect 8024 28364 8076 28416
rect 8852 28364 8904 28416
rect 9588 28407 9640 28416
rect 9588 28373 9597 28407
rect 9597 28373 9631 28407
rect 9631 28373 9640 28407
rect 9588 28364 9640 28373
rect 15292 28364 15344 28416
rect 18052 28407 18104 28416
rect 18052 28373 18061 28407
rect 18061 28373 18095 28407
rect 18095 28373 18104 28407
rect 18052 28364 18104 28373
rect 20352 28364 20404 28416
rect 35348 28509 35357 28543
rect 35357 28509 35391 28543
rect 35391 28509 35400 28543
rect 35348 28500 35400 28509
rect 36268 28500 36320 28552
rect 35164 28364 35216 28416
rect 15398 28262 15450 28314
rect 15462 28262 15514 28314
rect 15526 28262 15578 28314
rect 15590 28262 15642 28314
rect 15654 28262 15706 28314
rect 29846 28262 29898 28314
rect 29910 28262 29962 28314
rect 29974 28262 30026 28314
rect 30038 28262 30090 28314
rect 30102 28262 30154 28314
rect 44294 28262 44346 28314
rect 44358 28262 44410 28314
rect 44422 28262 44474 28314
rect 44486 28262 44538 28314
rect 44550 28262 44602 28314
rect 2320 28203 2372 28212
rect 2320 28169 2329 28203
rect 2329 28169 2363 28203
rect 2363 28169 2372 28203
rect 2320 28160 2372 28169
rect 6368 28203 6420 28212
rect 6368 28169 6377 28203
rect 6377 28169 6411 28203
rect 6411 28169 6420 28203
rect 6368 28160 6420 28169
rect 6460 28160 6512 28212
rect 18052 28160 18104 28212
rect 20628 28160 20680 28212
rect 37556 28160 37608 28212
rect 2780 28092 2832 28144
rect 4252 28092 4304 28144
rect 6276 28092 6328 28144
rect 5540 28024 5592 28076
rect 1860 27999 1912 28008
rect 1860 27965 1869 27999
rect 1869 27965 1903 27999
rect 1903 27965 1912 27999
rect 1860 27956 1912 27965
rect 2504 27956 2556 28008
rect 6644 27999 6696 28008
rect 6644 27965 6653 27999
rect 6653 27965 6687 27999
rect 6687 27965 6696 27999
rect 6644 27956 6696 27965
rect 7932 28092 7984 28144
rect 9128 28135 9180 28144
rect 9128 28101 9137 28135
rect 9137 28101 9171 28135
rect 9171 28101 9180 28135
rect 9128 28092 9180 28101
rect 18604 28092 18656 28144
rect 20352 28135 20404 28144
rect 20352 28101 20361 28135
rect 20361 28101 20395 28135
rect 20395 28101 20404 28135
rect 20352 28092 20404 28101
rect 7104 28024 7156 28076
rect 17776 27999 17828 28008
rect 8760 27888 8812 27940
rect 9680 27888 9732 27940
rect 17776 27965 17785 27999
rect 17785 27965 17819 27999
rect 17819 27965 17828 27999
rect 17776 27956 17828 27965
rect 34796 28024 34848 28076
rect 35348 28024 35400 28076
rect 36084 28067 36136 28076
rect 36084 28033 36093 28067
rect 36093 28033 36127 28067
rect 36127 28033 36136 28067
rect 36084 28024 36136 28033
rect 58072 28067 58124 28076
rect 58072 28033 58081 28067
rect 58081 28033 58115 28067
rect 58115 28033 58124 28067
rect 58072 28024 58124 28033
rect 35164 27999 35216 28008
rect 35164 27965 35173 27999
rect 35173 27965 35207 27999
rect 35207 27965 35216 27999
rect 35164 27956 35216 27965
rect 4344 27820 4396 27872
rect 16764 27863 16816 27872
rect 16764 27829 16773 27863
rect 16773 27829 16807 27863
rect 16807 27829 16816 27863
rect 16764 27820 16816 27829
rect 19340 27888 19392 27940
rect 57704 27888 57756 27940
rect 19616 27820 19668 27872
rect 34796 27820 34848 27872
rect 8174 27718 8226 27770
rect 8238 27718 8290 27770
rect 8302 27718 8354 27770
rect 8366 27718 8418 27770
rect 8430 27718 8482 27770
rect 22622 27718 22674 27770
rect 22686 27718 22738 27770
rect 22750 27718 22802 27770
rect 22814 27718 22866 27770
rect 22878 27718 22930 27770
rect 37070 27718 37122 27770
rect 37134 27718 37186 27770
rect 37198 27718 37250 27770
rect 37262 27718 37314 27770
rect 37326 27718 37378 27770
rect 51518 27718 51570 27770
rect 51582 27718 51634 27770
rect 51646 27718 51698 27770
rect 51710 27718 51762 27770
rect 51774 27718 51826 27770
rect 16764 27616 16816 27668
rect 17776 27616 17828 27668
rect 36084 27616 36136 27668
rect 40960 27616 41012 27668
rect 58072 27659 58124 27668
rect 58072 27625 58081 27659
rect 58081 27625 58115 27659
rect 58115 27625 58124 27659
rect 58072 27616 58124 27625
rect 4252 27591 4304 27600
rect 4252 27557 4261 27591
rect 4261 27557 4295 27591
rect 4295 27557 4304 27591
rect 4252 27548 4304 27557
rect 2872 27480 2924 27532
rect 4252 27412 4304 27464
rect 2504 27344 2556 27396
rect 3884 27344 3936 27396
rect 3700 27276 3752 27328
rect 4068 27276 4120 27328
rect 5448 27412 5500 27464
rect 9680 27523 9732 27532
rect 9680 27489 9689 27523
rect 9689 27489 9723 27523
rect 9723 27489 9732 27523
rect 9680 27480 9732 27489
rect 15292 27480 15344 27532
rect 19616 27523 19668 27532
rect 19616 27489 19625 27523
rect 19625 27489 19659 27523
rect 19659 27489 19668 27523
rect 19616 27480 19668 27489
rect 7472 27412 7524 27464
rect 8576 27412 8628 27464
rect 9404 27412 9456 27464
rect 14372 27412 14424 27464
rect 18236 27412 18288 27464
rect 7012 27344 7064 27396
rect 7932 27276 7984 27328
rect 8944 27319 8996 27328
rect 8944 27285 8953 27319
rect 8953 27285 8987 27319
rect 8987 27285 8996 27319
rect 8944 27276 8996 27285
rect 9588 27276 9640 27328
rect 10876 27276 10928 27328
rect 15752 27276 15804 27328
rect 18052 27344 18104 27396
rect 19432 27387 19484 27396
rect 19432 27353 19441 27387
rect 19441 27353 19475 27387
rect 19475 27353 19484 27387
rect 19432 27344 19484 27353
rect 45836 27344 45888 27396
rect 30288 27276 30340 27328
rect 35164 27276 35216 27328
rect 15398 27174 15450 27226
rect 15462 27174 15514 27226
rect 15526 27174 15578 27226
rect 15590 27174 15642 27226
rect 15654 27174 15706 27226
rect 29846 27174 29898 27226
rect 29910 27174 29962 27226
rect 29974 27174 30026 27226
rect 30038 27174 30090 27226
rect 30102 27174 30154 27226
rect 44294 27174 44346 27226
rect 44358 27174 44410 27226
rect 44422 27174 44474 27226
rect 44486 27174 44538 27226
rect 44550 27174 44602 27226
rect 2504 27072 2556 27124
rect 4160 27072 4212 27124
rect 5448 27115 5500 27124
rect 5448 27081 5457 27115
rect 5457 27081 5491 27115
rect 5491 27081 5500 27115
rect 5448 27072 5500 27081
rect 5540 27072 5592 27124
rect 8944 27072 8996 27124
rect 18052 27115 18104 27124
rect 18052 27081 18061 27115
rect 18061 27081 18095 27115
rect 18095 27081 18104 27115
rect 18052 27072 18104 27081
rect 3884 27047 3936 27056
rect 3884 27013 3893 27047
rect 3893 27013 3927 27047
rect 3927 27013 3936 27047
rect 3884 27004 3936 27013
rect 4068 27004 4120 27056
rect 3792 26936 3844 26988
rect 9956 27004 10008 27056
rect 15752 27004 15804 27056
rect 17684 27004 17736 27056
rect 7748 26936 7800 26988
rect 8024 26936 8076 26988
rect 14464 26979 14516 26988
rect 14464 26945 14473 26979
rect 14473 26945 14507 26979
rect 14507 26945 14516 26979
rect 14464 26936 14516 26945
rect 15292 26979 15344 26988
rect 15292 26945 15301 26979
rect 15301 26945 15335 26979
rect 15335 26945 15344 26979
rect 15292 26936 15344 26945
rect 17500 26936 17552 26988
rect 4068 26800 4120 26852
rect 7656 26868 7708 26920
rect 8944 26868 8996 26920
rect 14556 26911 14608 26920
rect 14556 26877 14565 26911
rect 14565 26877 14599 26911
rect 14599 26877 14608 26911
rect 14556 26868 14608 26877
rect 15936 26868 15988 26920
rect 23388 26936 23440 26988
rect 2412 26732 2464 26784
rect 4436 26732 4488 26784
rect 9864 26800 9916 26852
rect 13820 26800 13872 26852
rect 8576 26775 8628 26784
rect 8576 26741 8585 26775
rect 8585 26741 8619 26775
rect 8619 26741 8628 26775
rect 8576 26732 8628 26741
rect 12532 26732 12584 26784
rect 14188 26775 14240 26784
rect 14188 26741 14197 26775
rect 14197 26741 14231 26775
rect 14231 26741 14240 26775
rect 14188 26732 14240 26741
rect 20720 26800 20772 26852
rect 23020 26800 23072 26852
rect 17868 26732 17920 26784
rect 20076 26732 20128 26784
rect 24216 26775 24268 26784
rect 24216 26741 24225 26775
rect 24225 26741 24259 26775
rect 24259 26741 24268 26775
rect 24216 26732 24268 26741
rect 30288 26732 30340 26784
rect 8174 26630 8226 26682
rect 8238 26630 8290 26682
rect 8302 26630 8354 26682
rect 8366 26630 8418 26682
rect 8430 26630 8482 26682
rect 22622 26630 22674 26682
rect 22686 26630 22738 26682
rect 22750 26630 22802 26682
rect 22814 26630 22866 26682
rect 22878 26630 22930 26682
rect 37070 26630 37122 26682
rect 37134 26630 37186 26682
rect 37198 26630 37250 26682
rect 37262 26630 37314 26682
rect 37326 26630 37378 26682
rect 51518 26630 51570 26682
rect 51582 26630 51634 26682
rect 51646 26630 51698 26682
rect 51710 26630 51762 26682
rect 51774 26630 51826 26682
rect 3792 26571 3844 26580
rect 3792 26537 3801 26571
rect 3801 26537 3835 26571
rect 3835 26537 3844 26571
rect 3792 26528 3844 26537
rect 10876 26571 10928 26580
rect 10876 26537 10885 26571
rect 10885 26537 10919 26571
rect 10919 26537 10928 26571
rect 10876 26528 10928 26537
rect 5908 26460 5960 26512
rect 8024 26460 8076 26512
rect 12256 26460 12308 26512
rect 4068 26392 4120 26444
rect 5540 26435 5592 26444
rect 5540 26401 5549 26435
rect 5549 26401 5583 26435
rect 5583 26401 5592 26435
rect 5540 26392 5592 26401
rect 5724 26392 5776 26444
rect 6644 26435 6696 26444
rect 6644 26401 6653 26435
rect 6653 26401 6687 26435
rect 6687 26401 6696 26435
rect 6644 26392 6696 26401
rect 7932 26392 7984 26444
rect 2872 26324 2924 26376
rect 1676 26188 1728 26240
rect 3056 26188 3108 26240
rect 5816 26324 5868 26376
rect 5264 26299 5316 26308
rect 5264 26265 5273 26299
rect 5273 26265 5307 26299
rect 5307 26265 5316 26299
rect 5264 26256 5316 26265
rect 7748 26324 7800 26376
rect 9956 26392 10008 26444
rect 14648 26435 14700 26444
rect 14648 26401 14657 26435
rect 14657 26401 14691 26435
rect 14691 26401 14700 26435
rect 14648 26392 14700 26401
rect 15108 26435 15160 26444
rect 15108 26401 15117 26435
rect 15117 26401 15151 26435
rect 15151 26401 15160 26435
rect 15108 26392 15160 26401
rect 17224 26528 17276 26580
rect 17684 26528 17736 26580
rect 40776 26528 40828 26580
rect 18144 26503 18196 26512
rect 18144 26469 18153 26503
rect 18153 26469 18187 26503
rect 18187 26469 18196 26503
rect 18144 26460 18196 26469
rect 18972 26460 19024 26512
rect 23388 26460 23440 26512
rect 20352 26392 20404 26444
rect 24216 26392 24268 26444
rect 8944 26367 8996 26376
rect 8944 26333 8953 26367
rect 8953 26333 8987 26367
rect 8987 26333 8996 26367
rect 8944 26324 8996 26333
rect 9404 26324 9456 26376
rect 11060 26324 11112 26376
rect 13360 26367 13412 26376
rect 13360 26333 13369 26367
rect 13369 26333 13403 26367
rect 13403 26333 13412 26367
rect 13360 26324 13412 26333
rect 14464 26324 14516 26376
rect 15752 26367 15804 26376
rect 15752 26333 15761 26367
rect 15761 26333 15795 26367
rect 15795 26333 15804 26367
rect 15752 26324 15804 26333
rect 15844 26324 15896 26376
rect 17684 26367 17736 26376
rect 17684 26333 17693 26367
rect 17693 26333 17727 26367
rect 17727 26333 17736 26367
rect 17684 26324 17736 26333
rect 19616 26367 19668 26376
rect 19616 26333 19625 26367
rect 19625 26333 19659 26367
rect 19659 26333 19668 26367
rect 19616 26324 19668 26333
rect 20444 26367 20496 26376
rect 20444 26333 20453 26367
rect 20453 26333 20487 26367
rect 20487 26333 20496 26367
rect 20444 26324 20496 26333
rect 27344 26324 27396 26376
rect 37648 26324 37700 26376
rect 9220 26256 9272 26308
rect 9864 26256 9916 26308
rect 12532 26256 12584 26308
rect 13452 26299 13504 26308
rect 13452 26265 13461 26299
rect 13461 26265 13495 26299
rect 13495 26265 13504 26299
rect 13452 26256 13504 26265
rect 15016 26256 15068 26308
rect 22376 26299 22428 26308
rect 17040 26188 17092 26240
rect 20628 26231 20680 26240
rect 20628 26197 20637 26231
rect 20637 26197 20671 26231
rect 20671 26197 20680 26231
rect 20628 26188 20680 26197
rect 22376 26265 22385 26299
rect 22385 26265 22419 26299
rect 22419 26265 22428 26299
rect 22376 26256 22428 26265
rect 37556 26256 37608 26308
rect 23112 26188 23164 26240
rect 23848 26231 23900 26240
rect 23848 26197 23857 26231
rect 23857 26197 23891 26231
rect 23891 26197 23900 26231
rect 23848 26188 23900 26197
rect 15398 26086 15450 26138
rect 15462 26086 15514 26138
rect 15526 26086 15578 26138
rect 15590 26086 15642 26138
rect 15654 26086 15706 26138
rect 29846 26086 29898 26138
rect 29910 26086 29962 26138
rect 29974 26086 30026 26138
rect 30038 26086 30090 26138
rect 30102 26086 30154 26138
rect 44294 26086 44346 26138
rect 44358 26086 44410 26138
rect 44422 26086 44474 26138
rect 44486 26086 44538 26138
rect 44550 26086 44602 26138
rect 3976 25984 4028 26036
rect 7840 25984 7892 26036
rect 1676 25959 1728 25968
rect 1676 25925 1685 25959
rect 1685 25925 1719 25959
rect 1719 25925 1728 25959
rect 1676 25916 1728 25925
rect 9956 25916 10008 25968
rect 11060 25984 11112 26036
rect 15844 25984 15896 26036
rect 14188 25916 14240 25968
rect 15384 25916 15436 25968
rect 20444 25984 20496 26036
rect 22376 26027 22428 26036
rect 22376 25993 22385 26027
rect 22385 25993 22419 26027
rect 22419 25993 22428 26027
rect 22376 25984 22428 25993
rect 23388 25916 23440 25968
rect 30288 25959 30340 25968
rect 30288 25925 30297 25959
rect 30297 25925 30331 25959
rect 30331 25925 30340 25959
rect 30288 25916 30340 25925
rect 2780 25848 2832 25900
rect 3700 25891 3752 25900
rect 3700 25857 3709 25891
rect 3709 25857 3743 25891
rect 3743 25857 3752 25891
rect 3700 25848 3752 25857
rect 5264 25848 5316 25900
rect 5540 25848 5592 25900
rect 8576 25891 8628 25900
rect 7380 25780 7432 25832
rect 2872 25712 2924 25764
rect 3056 25644 3108 25696
rect 4804 25712 4856 25764
rect 8576 25857 8585 25891
rect 8585 25857 8619 25891
rect 8619 25857 8628 25891
rect 8576 25848 8628 25857
rect 9220 25891 9272 25900
rect 9220 25857 9229 25891
rect 9229 25857 9263 25891
rect 9263 25857 9272 25891
rect 9220 25848 9272 25857
rect 10968 25848 11020 25900
rect 13820 25891 13872 25900
rect 13820 25857 13829 25891
rect 13829 25857 13863 25891
rect 13863 25857 13872 25891
rect 13820 25848 13872 25857
rect 10876 25780 10928 25832
rect 11060 25780 11112 25832
rect 12256 25780 12308 25832
rect 14464 25780 14516 25832
rect 19616 25848 19668 25900
rect 20444 25891 20496 25900
rect 20444 25857 20453 25891
rect 20453 25857 20487 25891
rect 20487 25857 20496 25891
rect 20444 25848 20496 25857
rect 23848 25891 23900 25900
rect 17040 25823 17092 25832
rect 17040 25789 17049 25823
rect 17049 25789 17083 25823
rect 17083 25789 17092 25823
rect 17040 25780 17092 25789
rect 17868 25780 17920 25832
rect 18328 25823 18380 25832
rect 18328 25789 18337 25823
rect 18337 25789 18371 25823
rect 18371 25789 18380 25823
rect 18328 25780 18380 25789
rect 20352 25823 20404 25832
rect 20352 25789 20361 25823
rect 20361 25789 20395 25823
rect 20395 25789 20404 25823
rect 20352 25780 20404 25789
rect 20904 25780 20956 25832
rect 12532 25712 12584 25764
rect 13636 25712 13688 25764
rect 16672 25712 16724 25764
rect 17776 25712 17828 25764
rect 20812 25755 20864 25764
rect 20812 25721 20821 25755
rect 20821 25721 20855 25755
rect 20855 25721 20864 25755
rect 20812 25712 20864 25721
rect 21548 25712 21600 25764
rect 23848 25857 23857 25891
rect 23857 25857 23891 25891
rect 23891 25857 23900 25891
rect 23848 25848 23900 25857
rect 3608 25644 3660 25696
rect 3976 25644 4028 25696
rect 6828 25687 6880 25696
rect 6828 25653 6837 25687
rect 6837 25653 6871 25687
rect 6871 25653 6880 25687
rect 6828 25644 6880 25653
rect 7288 25644 7340 25696
rect 8668 25687 8720 25696
rect 8668 25653 8677 25687
rect 8677 25653 8711 25687
rect 8711 25653 8720 25687
rect 8668 25644 8720 25653
rect 12072 25687 12124 25696
rect 12072 25653 12081 25687
rect 12081 25653 12115 25687
rect 12115 25653 12124 25687
rect 12072 25644 12124 25653
rect 13544 25644 13596 25696
rect 19800 25644 19852 25696
rect 27436 25644 27488 25696
rect 28724 25848 28776 25900
rect 35992 25848 36044 25900
rect 30932 25687 30984 25696
rect 30932 25653 30941 25687
rect 30941 25653 30975 25687
rect 30975 25653 30984 25687
rect 30932 25644 30984 25653
rect 8174 25542 8226 25594
rect 8238 25542 8290 25594
rect 8302 25542 8354 25594
rect 8366 25542 8418 25594
rect 8430 25542 8482 25594
rect 22622 25542 22674 25594
rect 22686 25542 22738 25594
rect 22750 25542 22802 25594
rect 22814 25542 22866 25594
rect 22878 25542 22930 25594
rect 37070 25542 37122 25594
rect 37134 25542 37186 25594
rect 37198 25542 37250 25594
rect 37262 25542 37314 25594
rect 37326 25542 37378 25594
rect 51518 25542 51570 25594
rect 51582 25542 51634 25594
rect 51646 25542 51698 25594
rect 51710 25542 51762 25594
rect 51774 25542 51826 25594
rect 5540 25483 5592 25492
rect 5540 25449 5549 25483
rect 5549 25449 5583 25483
rect 5583 25449 5592 25483
rect 5540 25440 5592 25449
rect 9404 25440 9456 25492
rect 10876 25483 10928 25492
rect 10876 25449 10885 25483
rect 10885 25449 10919 25483
rect 10919 25449 10928 25483
rect 10876 25440 10928 25449
rect 9220 25372 9272 25424
rect 11152 25372 11204 25424
rect 7932 25347 7984 25356
rect 2412 25279 2464 25288
rect 1492 25143 1544 25152
rect 1492 25109 1501 25143
rect 1501 25109 1535 25143
rect 1535 25109 1544 25143
rect 1492 25100 1544 25109
rect 2412 25245 2421 25279
rect 2421 25245 2455 25279
rect 2455 25245 2464 25279
rect 2412 25236 2464 25245
rect 4344 25168 4396 25220
rect 7932 25313 7941 25347
rect 7941 25313 7975 25347
rect 7975 25313 7984 25347
rect 7932 25304 7984 25313
rect 11060 25304 11112 25356
rect 13268 25440 13320 25492
rect 18328 25440 18380 25492
rect 12164 25372 12216 25424
rect 14556 25372 14608 25424
rect 12348 25347 12400 25356
rect 12348 25313 12357 25347
rect 12357 25313 12391 25347
rect 12391 25313 12400 25347
rect 12348 25304 12400 25313
rect 12624 25347 12676 25356
rect 12624 25313 12633 25347
rect 12633 25313 12667 25347
rect 12667 25313 12676 25347
rect 12624 25304 12676 25313
rect 17592 25304 17644 25356
rect 7840 25279 7892 25288
rect 7840 25245 7849 25279
rect 7849 25245 7883 25279
rect 7883 25245 7892 25279
rect 7840 25236 7892 25245
rect 8944 25279 8996 25288
rect 8944 25245 8953 25279
rect 8953 25245 8987 25279
rect 8987 25245 8996 25279
rect 8944 25236 8996 25245
rect 9956 25279 10008 25288
rect 9956 25245 9965 25279
rect 9965 25245 9999 25279
rect 9999 25245 10008 25279
rect 9956 25236 10008 25245
rect 10968 25236 11020 25288
rect 3148 25143 3200 25152
rect 3148 25109 3157 25143
rect 3157 25109 3191 25143
rect 3191 25109 3200 25143
rect 3148 25100 3200 25109
rect 3516 25100 3568 25152
rect 6092 25143 6144 25152
rect 6092 25109 6101 25143
rect 6101 25109 6135 25143
rect 6135 25109 6144 25143
rect 6092 25100 6144 25109
rect 8024 25168 8076 25220
rect 12624 25168 12676 25220
rect 14648 25236 14700 25288
rect 15200 25236 15252 25288
rect 16028 25279 16080 25288
rect 16028 25245 16037 25279
rect 16037 25245 16071 25279
rect 16071 25245 16080 25279
rect 16028 25236 16080 25245
rect 17408 25236 17460 25288
rect 17776 25236 17828 25288
rect 18052 25415 18104 25424
rect 18052 25381 18061 25415
rect 18061 25381 18095 25415
rect 18095 25381 18104 25415
rect 18052 25372 18104 25381
rect 18328 25304 18380 25356
rect 19616 25304 19668 25356
rect 22284 25372 22336 25424
rect 20996 25304 21048 25356
rect 26332 25347 26384 25356
rect 26332 25313 26341 25347
rect 26341 25313 26375 25347
rect 26375 25313 26384 25347
rect 26332 25304 26384 25313
rect 19708 25236 19760 25288
rect 20352 25279 20404 25288
rect 20352 25245 20361 25279
rect 20361 25245 20395 25279
rect 20395 25245 20404 25279
rect 20352 25236 20404 25245
rect 20444 25236 20496 25288
rect 21456 25236 21508 25288
rect 21916 25236 21968 25288
rect 28724 25279 28776 25288
rect 28724 25245 28733 25279
rect 28733 25245 28767 25279
rect 28767 25245 28776 25279
rect 28724 25236 28776 25245
rect 29552 25279 29604 25288
rect 29552 25245 29561 25279
rect 29561 25245 29595 25279
rect 29595 25245 29604 25279
rect 29552 25236 29604 25245
rect 30932 25236 30984 25288
rect 31760 25279 31812 25288
rect 31760 25245 31769 25279
rect 31769 25245 31803 25279
rect 31803 25245 31812 25279
rect 31760 25236 31812 25245
rect 34980 25279 35032 25288
rect 34980 25245 34989 25279
rect 34989 25245 35023 25279
rect 35023 25245 35032 25279
rect 34980 25236 35032 25245
rect 7012 25100 7064 25152
rect 11428 25100 11480 25152
rect 12900 25100 12952 25152
rect 15936 25143 15988 25152
rect 15936 25109 15945 25143
rect 15945 25109 15979 25143
rect 15979 25109 15988 25143
rect 15936 25100 15988 25109
rect 18696 25100 18748 25152
rect 19524 25168 19576 25220
rect 20076 25168 20128 25220
rect 23940 25168 23992 25220
rect 26608 25211 26660 25220
rect 26608 25177 26617 25211
rect 26617 25177 26651 25211
rect 26651 25177 26660 25211
rect 26608 25168 26660 25177
rect 34520 25168 34572 25220
rect 21272 25100 21324 25152
rect 21456 25100 21508 25152
rect 22008 25100 22060 25152
rect 23204 25100 23256 25152
rect 28080 25143 28132 25152
rect 28080 25109 28089 25143
rect 28089 25109 28123 25143
rect 28123 25109 28132 25143
rect 28080 25100 28132 25109
rect 31300 25143 31352 25152
rect 31300 25109 31309 25143
rect 31309 25109 31343 25143
rect 31343 25109 31352 25143
rect 31300 25100 31352 25109
rect 15398 24998 15450 25050
rect 15462 24998 15514 25050
rect 15526 24998 15578 25050
rect 15590 24998 15642 25050
rect 15654 24998 15706 25050
rect 29846 24998 29898 25050
rect 29910 24998 29962 25050
rect 29974 24998 30026 25050
rect 30038 24998 30090 25050
rect 30102 24998 30154 25050
rect 44294 24998 44346 25050
rect 44358 24998 44410 25050
rect 44422 24998 44474 25050
rect 44486 24998 44538 25050
rect 44550 24998 44602 25050
rect 4344 24896 4396 24948
rect 3700 24803 3752 24812
rect 3700 24769 3709 24803
rect 3709 24769 3743 24803
rect 3743 24769 3752 24803
rect 3700 24760 3752 24769
rect 4804 24803 4856 24812
rect 4804 24769 4813 24803
rect 4813 24769 4847 24803
rect 4847 24769 4856 24803
rect 4804 24760 4856 24769
rect 3608 24735 3660 24744
rect 3608 24701 3617 24735
rect 3617 24701 3651 24735
rect 3651 24701 3660 24735
rect 3608 24692 3660 24701
rect 6092 24828 6144 24880
rect 5632 24803 5684 24812
rect 5632 24769 5641 24803
rect 5641 24769 5675 24803
rect 5675 24769 5684 24803
rect 5632 24760 5684 24769
rect 7288 24828 7340 24880
rect 9680 24828 9732 24880
rect 12624 24871 12676 24880
rect 12624 24837 12633 24871
rect 12633 24837 12667 24871
rect 12667 24837 12676 24871
rect 12624 24828 12676 24837
rect 8668 24760 8720 24812
rect 10968 24760 11020 24812
rect 12256 24760 12308 24812
rect 12900 24760 12952 24812
rect 16028 24896 16080 24948
rect 21824 24896 21876 24948
rect 22008 24896 22060 24948
rect 22376 24896 22428 24948
rect 26608 24896 26660 24948
rect 19800 24828 19852 24880
rect 29552 24828 29604 24880
rect 3056 24667 3108 24676
rect 3056 24633 3065 24667
rect 3065 24633 3099 24667
rect 3099 24633 3108 24667
rect 3056 24624 3108 24633
rect 6552 24624 6604 24676
rect 1952 24599 2004 24608
rect 1952 24565 1961 24599
rect 1961 24565 1995 24599
rect 1995 24565 2004 24599
rect 1952 24556 2004 24565
rect 2228 24556 2280 24608
rect 4896 24556 4948 24608
rect 8760 24692 8812 24744
rect 9220 24735 9272 24744
rect 9220 24701 9229 24735
rect 9229 24701 9263 24735
rect 9263 24701 9272 24735
rect 9220 24692 9272 24701
rect 13728 24624 13780 24676
rect 7380 24556 7432 24608
rect 9680 24556 9732 24608
rect 10692 24599 10744 24608
rect 10692 24565 10701 24599
rect 10701 24565 10735 24599
rect 10735 24565 10744 24599
rect 10692 24556 10744 24565
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 14924 24692 14976 24744
rect 17316 24760 17368 24812
rect 18328 24760 18380 24812
rect 18788 24760 18840 24812
rect 19156 24760 19208 24812
rect 15200 24692 15252 24744
rect 17040 24692 17092 24744
rect 17592 24735 17644 24744
rect 17592 24701 17601 24735
rect 17601 24701 17635 24735
rect 17635 24701 17644 24735
rect 17592 24692 17644 24701
rect 21272 24760 21324 24812
rect 22008 24803 22060 24812
rect 19616 24735 19668 24744
rect 19616 24701 19625 24735
rect 19625 24701 19659 24735
rect 19659 24701 19668 24735
rect 19616 24692 19668 24701
rect 20628 24692 20680 24744
rect 18512 24624 18564 24676
rect 21088 24735 21140 24744
rect 21088 24701 21097 24735
rect 21097 24701 21131 24735
rect 21131 24701 21140 24735
rect 22008 24769 22017 24803
rect 22017 24769 22051 24803
rect 22051 24769 22060 24803
rect 22008 24760 22060 24769
rect 24492 24803 24544 24812
rect 24492 24769 24501 24803
rect 24501 24769 24535 24803
rect 24535 24769 24544 24803
rect 24492 24760 24544 24769
rect 25044 24760 25096 24812
rect 26424 24803 26476 24812
rect 26424 24769 26433 24803
rect 26433 24769 26467 24803
rect 26467 24769 26476 24803
rect 26424 24760 26476 24769
rect 28080 24760 28132 24812
rect 29000 24803 29052 24812
rect 21088 24692 21140 24701
rect 21916 24692 21968 24744
rect 23388 24692 23440 24744
rect 25320 24735 25372 24744
rect 25320 24701 25329 24735
rect 25329 24701 25363 24735
rect 25363 24701 25372 24735
rect 25320 24692 25372 24701
rect 15844 24556 15896 24608
rect 16120 24556 16172 24608
rect 18144 24599 18196 24608
rect 18144 24565 18153 24599
rect 18153 24565 18187 24599
rect 18187 24565 18196 24599
rect 18144 24556 18196 24565
rect 19892 24599 19944 24608
rect 19892 24565 19901 24599
rect 19901 24565 19935 24599
rect 19935 24565 19944 24599
rect 19892 24556 19944 24565
rect 20536 24599 20588 24608
rect 20536 24565 20545 24599
rect 20545 24565 20579 24599
rect 20579 24565 20588 24599
rect 20536 24556 20588 24565
rect 22192 24624 22244 24676
rect 29000 24769 29009 24803
rect 29009 24769 29043 24803
rect 29043 24769 29052 24803
rect 29000 24760 29052 24769
rect 31760 24760 31812 24812
rect 35992 24803 36044 24812
rect 35992 24769 36001 24803
rect 36001 24769 36035 24803
rect 36035 24769 36044 24803
rect 35992 24760 36044 24769
rect 39028 24760 39080 24812
rect 31300 24692 31352 24744
rect 33416 24692 33468 24744
rect 33600 24735 33652 24744
rect 33600 24701 33609 24735
rect 33609 24701 33643 24735
rect 33643 24701 33652 24735
rect 33600 24692 33652 24701
rect 34520 24692 34572 24744
rect 37372 24735 37424 24744
rect 37372 24701 37381 24735
rect 37381 24701 37415 24735
rect 37415 24701 37424 24735
rect 37372 24692 37424 24701
rect 39948 24692 40000 24744
rect 31852 24624 31904 24676
rect 21640 24556 21692 24608
rect 21916 24599 21968 24608
rect 21916 24565 21925 24599
rect 21925 24565 21959 24599
rect 21959 24565 21968 24599
rect 21916 24556 21968 24565
rect 23756 24556 23808 24608
rect 23848 24599 23900 24608
rect 23848 24565 23857 24599
rect 23857 24565 23891 24599
rect 23891 24565 23900 24599
rect 23848 24556 23900 24565
rect 26792 24556 26844 24608
rect 28356 24599 28408 24608
rect 28356 24565 28365 24599
rect 28365 24565 28399 24599
rect 28399 24565 28408 24599
rect 28356 24556 28408 24565
rect 29736 24556 29788 24608
rect 30012 24599 30064 24608
rect 30012 24565 30021 24599
rect 30021 24565 30055 24599
rect 30055 24565 30064 24599
rect 30012 24556 30064 24565
rect 35348 24599 35400 24608
rect 35348 24565 35357 24599
rect 35357 24565 35391 24599
rect 35391 24565 35400 24599
rect 35348 24556 35400 24565
rect 39120 24599 39172 24608
rect 39120 24565 39129 24599
rect 39129 24565 39163 24599
rect 39163 24565 39172 24599
rect 39120 24556 39172 24565
rect 8174 24454 8226 24506
rect 8238 24454 8290 24506
rect 8302 24454 8354 24506
rect 8366 24454 8418 24506
rect 8430 24454 8482 24506
rect 22622 24454 22674 24506
rect 22686 24454 22738 24506
rect 22750 24454 22802 24506
rect 22814 24454 22866 24506
rect 22878 24454 22930 24506
rect 37070 24454 37122 24506
rect 37134 24454 37186 24506
rect 37198 24454 37250 24506
rect 37262 24454 37314 24506
rect 37326 24454 37378 24506
rect 51518 24454 51570 24506
rect 51582 24454 51634 24506
rect 51646 24454 51698 24506
rect 51710 24454 51762 24506
rect 51774 24454 51826 24506
rect 3148 24191 3200 24200
rect 3148 24157 3157 24191
rect 3157 24157 3191 24191
rect 3191 24157 3200 24191
rect 4160 24216 4212 24268
rect 3148 24148 3200 24157
rect 5724 24284 5776 24336
rect 7656 24327 7708 24336
rect 7656 24293 7665 24327
rect 7665 24293 7699 24327
rect 7699 24293 7708 24327
rect 7656 24284 7708 24293
rect 8116 24259 8168 24268
rect 8116 24225 8125 24259
rect 8125 24225 8159 24259
rect 8159 24225 8168 24259
rect 8116 24216 8168 24225
rect 9956 24352 10008 24404
rect 11704 24352 11756 24404
rect 13360 24352 13412 24404
rect 14464 24352 14516 24404
rect 14924 24352 14976 24404
rect 8760 24284 8812 24336
rect 5540 24191 5592 24200
rect 2872 24123 2924 24132
rect 2044 24012 2096 24064
rect 2872 24089 2881 24123
rect 2881 24089 2915 24123
rect 2915 24089 2924 24123
rect 2872 24080 2924 24089
rect 3332 24080 3384 24132
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 5632 24148 5684 24200
rect 7564 24148 7616 24200
rect 7840 24148 7892 24200
rect 4896 24080 4948 24132
rect 2780 24012 2832 24064
rect 3516 24012 3568 24064
rect 3792 24055 3844 24064
rect 3792 24021 3801 24055
rect 3801 24021 3835 24055
rect 3835 24021 3844 24055
rect 3792 24012 3844 24021
rect 10692 24216 10744 24268
rect 13268 24216 13320 24268
rect 13360 24216 13412 24268
rect 9680 24191 9732 24200
rect 9680 24157 9689 24191
rect 9689 24157 9723 24191
rect 9723 24157 9732 24191
rect 9680 24148 9732 24157
rect 12256 24148 12308 24200
rect 14648 24191 14700 24200
rect 14648 24157 14657 24191
rect 14657 24157 14691 24191
rect 14691 24157 14700 24191
rect 14648 24148 14700 24157
rect 15292 24191 15344 24200
rect 15292 24157 15301 24191
rect 15301 24157 15335 24191
rect 15335 24157 15344 24191
rect 15292 24148 15344 24157
rect 10968 24080 11020 24132
rect 15200 24080 15252 24132
rect 17592 24352 17644 24404
rect 23388 24352 23440 24404
rect 22008 24284 22060 24336
rect 17040 24148 17092 24200
rect 18328 24191 18380 24200
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 19064 24216 19116 24268
rect 19616 24216 19668 24268
rect 21824 24216 21876 24268
rect 22284 24216 22336 24268
rect 21364 24191 21416 24200
rect 21364 24157 21373 24191
rect 21373 24157 21407 24191
rect 21407 24157 21416 24191
rect 21364 24148 21416 24157
rect 22100 24148 22152 24200
rect 23204 24148 23256 24200
rect 25136 24284 25188 24336
rect 26424 24352 26476 24404
rect 27988 24352 28040 24404
rect 29000 24395 29052 24404
rect 29000 24361 29009 24395
rect 29009 24361 29043 24395
rect 29043 24361 29052 24395
rect 29000 24352 29052 24361
rect 30012 24352 30064 24404
rect 31760 24352 31812 24404
rect 33416 24352 33468 24404
rect 24124 24216 24176 24268
rect 26424 24216 26476 24268
rect 28724 24216 28776 24268
rect 34980 24352 35032 24404
rect 35992 24352 36044 24404
rect 37740 24352 37792 24404
rect 38568 24352 38620 24404
rect 39028 24395 39080 24404
rect 39028 24361 39037 24395
rect 39037 24361 39071 24395
rect 39071 24361 39080 24395
rect 39028 24352 39080 24361
rect 39948 24395 40000 24404
rect 39948 24361 39957 24395
rect 39957 24361 39991 24395
rect 39991 24361 40000 24395
rect 39948 24352 40000 24361
rect 40684 24284 40736 24336
rect 23756 24148 23808 24200
rect 26516 24191 26568 24200
rect 26516 24157 26525 24191
rect 26525 24157 26559 24191
rect 26559 24157 26568 24191
rect 26516 24148 26568 24157
rect 18144 24080 18196 24132
rect 23848 24080 23900 24132
rect 26792 24123 26844 24132
rect 20444 24012 20496 24064
rect 20996 24012 21048 24064
rect 22468 24055 22520 24064
rect 22468 24021 22477 24055
rect 22477 24021 22511 24055
rect 22511 24021 22520 24055
rect 22468 24012 22520 24021
rect 24768 24012 24820 24064
rect 25136 24012 25188 24064
rect 26240 24012 26292 24064
rect 26792 24089 26801 24123
rect 26801 24089 26835 24123
rect 26835 24089 26844 24123
rect 26792 24080 26844 24089
rect 28356 24080 28408 24132
rect 29552 24148 29604 24200
rect 31208 24080 31260 24132
rect 29460 24012 29512 24064
rect 31760 24012 31812 24064
rect 34980 24148 35032 24200
rect 35348 24148 35400 24200
rect 39120 24216 39172 24268
rect 38568 24148 38620 24200
rect 39856 24191 39908 24200
rect 39856 24157 39865 24191
rect 39865 24157 39899 24191
rect 39899 24157 39908 24191
rect 39856 24148 39908 24157
rect 33968 24080 34020 24132
rect 48320 24080 48372 24132
rect 37556 24012 37608 24064
rect 47584 24055 47636 24064
rect 47584 24021 47593 24055
rect 47593 24021 47627 24055
rect 47627 24021 47636 24055
rect 47584 24012 47636 24021
rect 15398 23910 15450 23962
rect 15462 23910 15514 23962
rect 15526 23910 15578 23962
rect 15590 23910 15642 23962
rect 15654 23910 15706 23962
rect 29846 23910 29898 23962
rect 29910 23910 29962 23962
rect 29974 23910 30026 23962
rect 30038 23910 30090 23962
rect 30102 23910 30154 23962
rect 44294 23910 44346 23962
rect 44358 23910 44410 23962
rect 44422 23910 44474 23962
rect 44486 23910 44538 23962
rect 44550 23910 44602 23962
rect 2964 23740 3016 23792
rect 5816 23808 5868 23860
rect 9036 23808 9088 23860
rect 9312 23808 9364 23860
rect 15200 23851 15252 23860
rect 15200 23817 15209 23851
rect 15209 23817 15243 23851
rect 15243 23817 15252 23851
rect 15200 23808 15252 23817
rect 22468 23808 22520 23860
rect 25136 23808 25188 23860
rect 31208 23808 31260 23860
rect 6092 23740 6144 23792
rect 13176 23740 13228 23792
rect 14648 23740 14700 23792
rect 24584 23783 24636 23792
rect 2044 23715 2096 23724
rect 2044 23681 2053 23715
rect 2053 23681 2087 23715
rect 2087 23681 2096 23715
rect 2044 23672 2096 23681
rect 3056 23715 3108 23724
rect 3056 23681 3065 23715
rect 3065 23681 3099 23715
rect 3099 23681 3108 23715
rect 3056 23672 3108 23681
rect 3332 23715 3384 23724
rect 3332 23681 3341 23715
rect 3341 23681 3375 23715
rect 3375 23681 3384 23715
rect 3332 23672 3384 23681
rect 3976 23715 4028 23724
rect 3976 23681 3985 23715
rect 3985 23681 4019 23715
rect 4019 23681 4028 23715
rect 3976 23672 4028 23681
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 3240 23536 3292 23588
rect 6000 23604 6052 23656
rect 6644 23672 6696 23724
rect 8576 23604 8628 23656
rect 9128 23604 9180 23656
rect 13452 23715 13504 23724
rect 13452 23681 13461 23715
rect 13461 23681 13495 23715
rect 13495 23681 13504 23715
rect 13912 23715 13964 23724
rect 13452 23672 13504 23681
rect 13912 23681 13921 23715
rect 13921 23681 13955 23715
rect 13955 23681 13964 23715
rect 13912 23672 13964 23681
rect 24584 23749 24593 23783
rect 24593 23749 24627 23783
rect 24627 23749 24636 23783
rect 24584 23740 24636 23749
rect 13084 23604 13136 23656
rect 16120 23604 16172 23656
rect 6368 23536 6420 23588
rect 7840 23536 7892 23588
rect 13452 23536 13504 23588
rect 13728 23536 13780 23588
rect 2228 23511 2280 23520
rect 2228 23477 2237 23511
rect 2237 23477 2271 23511
rect 2271 23477 2280 23511
rect 2228 23468 2280 23477
rect 4160 23468 4212 23520
rect 5632 23511 5684 23520
rect 5632 23477 5641 23511
rect 5641 23477 5675 23511
rect 5675 23477 5684 23511
rect 5632 23468 5684 23477
rect 5816 23511 5868 23520
rect 5816 23477 5825 23511
rect 5825 23477 5859 23511
rect 5859 23477 5868 23511
rect 5816 23468 5868 23477
rect 8024 23468 8076 23520
rect 9680 23511 9732 23520
rect 9680 23477 9689 23511
rect 9689 23477 9723 23511
rect 9723 23477 9732 23511
rect 9680 23468 9732 23477
rect 18328 23672 18380 23724
rect 17316 23604 17368 23656
rect 19616 23604 19668 23656
rect 19984 23647 20036 23656
rect 19984 23613 19993 23647
rect 19993 23613 20027 23647
rect 20027 23613 20036 23647
rect 19984 23604 20036 23613
rect 21180 23672 21232 23724
rect 21916 23672 21968 23724
rect 22008 23672 22060 23724
rect 24400 23672 24452 23724
rect 26424 23672 26476 23724
rect 26976 23672 27028 23724
rect 27988 23715 28040 23724
rect 27988 23681 27997 23715
rect 27997 23681 28031 23715
rect 28031 23681 28040 23715
rect 27988 23672 28040 23681
rect 47584 23808 47636 23860
rect 33876 23740 33928 23792
rect 35992 23740 36044 23792
rect 37556 23783 37608 23792
rect 37556 23749 37565 23783
rect 37565 23749 37599 23783
rect 37599 23749 37608 23783
rect 37556 23740 37608 23749
rect 40684 23740 40736 23792
rect 29552 23715 29604 23724
rect 29552 23681 29561 23715
rect 29561 23681 29595 23715
rect 29595 23681 29604 23715
rect 29552 23672 29604 23681
rect 29828 23672 29880 23724
rect 31852 23672 31904 23724
rect 32680 23672 32732 23724
rect 38660 23672 38712 23724
rect 39120 23672 39172 23724
rect 56600 23672 56652 23724
rect 21456 23604 21508 23656
rect 20260 23536 20312 23588
rect 24492 23604 24544 23656
rect 25504 23604 25556 23656
rect 28080 23647 28132 23656
rect 28080 23613 28089 23647
rect 28089 23613 28123 23647
rect 28123 23613 28132 23647
rect 28080 23604 28132 23613
rect 29276 23647 29328 23656
rect 29276 23613 29285 23647
rect 29285 23613 29319 23647
rect 29319 23613 29328 23647
rect 29276 23604 29328 23613
rect 29460 23647 29512 23656
rect 29460 23613 29469 23647
rect 29469 23613 29503 23647
rect 29503 23613 29512 23647
rect 29460 23604 29512 23613
rect 29644 23647 29696 23656
rect 29644 23613 29653 23647
rect 29653 23613 29687 23647
rect 29687 23613 29696 23647
rect 29644 23604 29696 23613
rect 23388 23536 23440 23588
rect 26608 23536 26660 23588
rect 27528 23536 27580 23588
rect 36544 23604 36596 23656
rect 39856 23604 39908 23656
rect 42708 23604 42760 23656
rect 47492 23604 47544 23656
rect 48596 23647 48648 23656
rect 48596 23613 48605 23647
rect 48605 23613 48639 23647
rect 48639 23613 48648 23647
rect 48596 23604 48648 23613
rect 19156 23511 19208 23520
rect 19156 23477 19165 23511
rect 19165 23477 19199 23511
rect 19199 23477 19208 23511
rect 19156 23468 19208 23477
rect 21824 23468 21876 23520
rect 23572 23468 23624 23520
rect 24124 23468 24176 23520
rect 24676 23468 24728 23520
rect 26056 23468 26108 23520
rect 28724 23468 28776 23520
rect 32128 23468 32180 23520
rect 35900 23468 35952 23520
rect 57888 23468 57940 23520
rect 8174 23366 8226 23418
rect 8238 23366 8290 23418
rect 8302 23366 8354 23418
rect 8366 23366 8418 23418
rect 8430 23366 8482 23418
rect 22622 23366 22674 23418
rect 22686 23366 22738 23418
rect 22750 23366 22802 23418
rect 22814 23366 22866 23418
rect 22878 23366 22930 23418
rect 37070 23366 37122 23418
rect 37134 23366 37186 23418
rect 37198 23366 37250 23418
rect 37262 23366 37314 23418
rect 37326 23366 37378 23418
rect 51518 23366 51570 23418
rect 51582 23366 51634 23418
rect 51646 23366 51698 23418
rect 51710 23366 51762 23418
rect 51774 23366 51826 23418
rect 3976 23264 4028 23316
rect 2872 23196 2924 23248
rect 3240 23128 3292 23180
rect 4528 23128 4580 23180
rect 6552 23171 6604 23180
rect 6552 23137 6561 23171
rect 6561 23137 6595 23171
rect 6595 23137 6604 23171
rect 6552 23128 6604 23137
rect 7564 23264 7616 23316
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 15384 23264 15436 23316
rect 18052 23264 18104 23316
rect 18328 23307 18380 23316
rect 18328 23273 18337 23307
rect 18337 23273 18371 23307
rect 18371 23273 18380 23307
rect 18328 23264 18380 23273
rect 18604 23264 18656 23316
rect 19524 23264 19576 23316
rect 22192 23307 22244 23316
rect 11152 23128 11204 23180
rect 2044 23103 2096 23112
rect 2044 23069 2053 23103
rect 2053 23069 2087 23103
rect 2087 23069 2096 23103
rect 2044 23060 2096 23069
rect 2228 23060 2280 23112
rect 3884 23103 3936 23112
rect 2780 22924 2832 22976
rect 3884 23069 3893 23103
rect 3893 23069 3927 23103
rect 3927 23069 3936 23103
rect 3884 23060 3936 23069
rect 9680 23060 9732 23112
rect 11060 23060 11112 23112
rect 13636 23128 13688 23180
rect 17040 23196 17092 23248
rect 17224 23239 17276 23248
rect 17224 23205 17233 23239
rect 17233 23205 17267 23239
rect 17267 23205 17276 23239
rect 17224 23196 17276 23205
rect 11796 23103 11848 23112
rect 11796 23069 11805 23103
rect 11805 23069 11839 23103
rect 11839 23069 11848 23103
rect 11796 23060 11848 23069
rect 13176 23060 13228 23112
rect 4620 22992 4672 23044
rect 6828 23035 6880 23044
rect 5540 22924 5592 22976
rect 6828 23001 6837 23035
rect 6837 23001 6871 23035
rect 6871 23001 6880 23035
rect 6828 22992 6880 23001
rect 7564 22992 7616 23044
rect 10140 22924 10192 22976
rect 12164 22992 12216 23044
rect 15936 23128 15988 23180
rect 19432 23196 19484 23248
rect 22192 23273 22201 23307
rect 22201 23273 22235 23307
rect 22235 23273 22244 23307
rect 27436 23307 27488 23316
rect 22192 23264 22244 23273
rect 18880 23128 18932 23180
rect 19524 23128 19576 23180
rect 20076 23128 20128 23180
rect 20996 23171 21048 23180
rect 20996 23137 21005 23171
rect 21005 23137 21039 23171
rect 21039 23137 21048 23171
rect 20996 23128 21048 23137
rect 22376 23196 22428 23248
rect 23940 23196 23992 23248
rect 23572 23128 23624 23180
rect 17408 23103 17460 23112
rect 15016 22992 15068 23044
rect 16212 22992 16264 23044
rect 16304 22924 16356 22976
rect 16764 22924 16816 22976
rect 17408 23069 17417 23103
rect 17417 23069 17451 23103
rect 17451 23069 17460 23103
rect 17408 23060 17460 23069
rect 18972 23060 19024 23112
rect 19984 23060 20036 23112
rect 20444 23060 20496 23112
rect 21180 23060 21232 23112
rect 21640 23060 21692 23112
rect 17960 22992 18012 23044
rect 18052 23035 18104 23044
rect 18052 23001 18061 23035
rect 18061 23001 18095 23035
rect 18095 23001 18104 23035
rect 18052 22992 18104 23001
rect 19248 22992 19300 23044
rect 19708 23035 19760 23044
rect 19708 23001 19717 23035
rect 19717 23001 19751 23035
rect 19751 23001 19760 23035
rect 19708 22992 19760 23001
rect 21364 23035 21416 23044
rect 21364 23001 21373 23035
rect 21373 23001 21407 23035
rect 21407 23001 21416 23035
rect 21364 22992 21416 23001
rect 23480 23035 23532 23044
rect 20536 22924 20588 22976
rect 23480 23001 23489 23035
rect 23489 23001 23523 23035
rect 23523 23001 23532 23035
rect 23480 22992 23532 23001
rect 24584 23103 24636 23112
rect 24584 23069 24593 23103
rect 24593 23069 24627 23103
rect 24627 23069 24636 23103
rect 24584 23060 24636 23069
rect 23572 22924 23624 22976
rect 24492 22992 24544 23044
rect 25596 23128 25648 23180
rect 27436 23273 27445 23307
rect 27445 23273 27479 23307
rect 27479 23273 27488 23307
rect 27436 23264 27488 23273
rect 27620 23264 27672 23316
rect 33968 23307 34020 23316
rect 33968 23273 33977 23307
rect 33977 23273 34011 23307
rect 34011 23273 34020 23307
rect 33968 23264 34020 23273
rect 35992 23307 36044 23316
rect 35992 23273 36001 23307
rect 36001 23273 36035 23307
rect 36035 23273 36044 23307
rect 35992 23264 36044 23273
rect 38660 23264 38712 23316
rect 28080 23239 28132 23248
rect 28080 23205 28089 23239
rect 28089 23205 28123 23239
rect 28123 23205 28132 23239
rect 28080 23196 28132 23205
rect 28632 23171 28684 23180
rect 28632 23137 28641 23171
rect 28641 23137 28675 23171
rect 28675 23137 28684 23171
rect 28632 23128 28684 23137
rect 31852 23128 31904 23180
rect 24952 23060 25004 23112
rect 25688 23103 25740 23112
rect 25688 23069 25697 23103
rect 25697 23069 25731 23103
rect 25731 23069 25740 23103
rect 25688 23060 25740 23069
rect 25780 23103 25832 23112
rect 25780 23069 25789 23103
rect 25789 23069 25823 23103
rect 25823 23069 25832 23103
rect 25780 23060 25832 23069
rect 26424 23060 26476 23112
rect 26608 23103 26660 23112
rect 26608 23069 26617 23103
rect 26617 23069 26651 23103
rect 26651 23069 26660 23103
rect 26884 23103 26936 23112
rect 26608 23060 26660 23069
rect 26884 23069 26893 23103
rect 26893 23069 26927 23103
rect 26927 23069 26936 23103
rect 26884 23060 26936 23069
rect 26976 23103 27028 23112
rect 26976 23069 26985 23103
rect 26985 23069 27019 23103
rect 27019 23069 27028 23103
rect 26976 23060 27028 23069
rect 28172 23060 28224 23112
rect 29000 23060 29052 23112
rect 36268 23128 36320 23180
rect 42524 23171 42576 23180
rect 35440 23103 35492 23112
rect 27988 22992 28040 23044
rect 35440 23069 35449 23103
rect 35449 23069 35483 23103
rect 35483 23069 35492 23103
rect 35440 23060 35492 23069
rect 31392 23035 31444 23044
rect 25136 22924 25188 22976
rect 25780 22924 25832 22976
rect 31392 23001 31401 23035
rect 31401 23001 31435 23035
rect 31435 23001 31444 23035
rect 31392 22992 31444 23001
rect 32128 22992 32180 23044
rect 32680 22992 32732 23044
rect 36360 23060 36412 23112
rect 42524 23137 42533 23171
rect 42533 23137 42567 23171
rect 42567 23137 42576 23171
rect 42524 23128 42576 23137
rect 42708 23128 42760 23180
rect 47584 23128 47636 23180
rect 48596 23171 48648 23180
rect 48596 23137 48605 23171
rect 48605 23137 48639 23171
rect 48639 23137 48648 23171
rect 48596 23128 48648 23137
rect 38384 23060 38436 23112
rect 43352 23103 43404 23112
rect 43352 23069 43361 23103
rect 43361 23069 43395 23103
rect 43395 23069 43404 23103
rect 47768 23103 47820 23112
rect 43352 23060 43404 23069
rect 47768 23069 47777 23103
rect 47777 23069 47811 23103
rect 47811 23069 47820 23103
rect 47768 23060 47820 23069
rect 28540 22967 28592 22976
rect 28540 22933 28549 22967
rect 28549 22933 28583 22967
rect 28583 22933 28592 22967
rect 28540 22924 28592 22933
rect 28816 22967 28868 22976
rect 28816 22933 28825 22967
rect 28825 22933 28859 22967
rect 28859 22933 28868 22967
rect 28816 22924 28868 22933
rect 32864 22967 32916 22976
rect 32864 22933 32873 22967
rect 32873 22933 32907 22967
rect 32907 22933 32916 22967
rect 32864 22924 32916 22933
rect 35072 22924 35124 22976
rect 46572 22924 46624 22976
rect 47400 22924 47452 22976
rect 15398 22822 15450 22874
rect 15462 22822 15514 22874
rect 15526 22822 15578 22874
rect 15590 22822 15642 22874
rect 15654 22822 15706 22874
rect 29846 22822 29898 22874
rect 29910 22822 29962 22874
rect 29974 22822 30026 22874
rect 30038 22822 30090 22874
rect 30102 22822 30154 22874
rect 44294 22822 44346 22874
rect 44358 22822 44410 22874
rect 44422 22822 44474 22874
rect 44486 22822 44538 22874
rect 44550 22822 44602 22874
rect 6644 22720 6696 22772
rect 6736 22720 6788 22772
rect 6920 22720 6972 22772
rect 7748 22720 7800 22772
rect 8024 22720 8076 22772
rect 3056 22652 3108 22704
rect 4712 22584 4764 22636
rect 7012 22652 7064 22704
rect 7656 22652 7708 22704
rect 6368 22584 6420 22636
rect 9772 22652 9824 22704
rect 13268 22720 13320 22772
rect 13728 22720 13780 22772
rect 14924 22720 14976 22772
rect 11060 22652 11112 22704
rect 6644 22516 6696 22568
rect 7104 22516 7156 22568
rect 7748 22516 7800 22568
rect 12532 22625 12584 22636
rect 12532 22591 12541 22625
rect 12541 22591 12575 22625
rect 12575 22591 12584 22625
rect 13176 22627 13228 22636
rect 12532 22584 12584 22591
rect 13176 22593 13185 22627
rect 13185 22593 13219 22627
rect 13219 22593 13228 22627
rect 13176 22584 13228 22593
rect 14096 22652 14148 22704
rect 17040 22720 17092 22772
rect 17316 22720 17368 22772
rect 20904 22720 20956 22772
rect 21272 22720 21324 22772
rect 16028 22584 16080 22636
rect 16304 22584 16356 22636
rect 17408 22584 17460 22636
rect 17776 22584 17828 22636
rect 23480 22652 23532 22704
rect 24216 22720 24268 22772
rect 24584 22720 24636 22772
rect 24676 22720 24728 22772
rect 25320 22763 25372 22772
rect 20720 22584 20772 22636
rect 2964 22448 3016 22500
rect 4988 22423 5040 22432
rect 4988 22389 4997 22423
rect 4997 22389 5031 22423
rect 5031 22389 5040 22423
rect 4988 22380 5040 22389
rect 5816 22380 5868 22432
rect 6000 22380 6052 22432
rect 15292 22516 15344 22568
rect 16580 22516 16632 22568
rect 11152 22448 11204 22500
rect 12440 22423 12492 22432
rect 12440 22389 12449 22423
rect 12449 22389 12483 22423
rect 12483 22389 12492 22423
rect 17132 22448 17184 22500
rect 18420 22491 18472 22500
rect 18420 22457 18429 22491
rect 18429 22457 18463 22491
rect 18463 22457 18472 22491
rect 18420 22448 18472 22457
rect 22284 22584 22336 22636
rect 21824 22559 21876 22568
rect 21824 22525 21833 22559
rect 21833 22525 21867 22559
rect 21867 22525 21876 22559
rect 21824 22516 21876 22525
rect 23664 22584 23716 22636
rect 23848 22627 23900 22636
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 23848 22584 23900 22593
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24676 22584 24728 22636
rect 25320 22729 25329 22763
rect 25329 22729 25363 22763
rect 25363 22729 25372 22763
rect 25320 22720 25372 22729
rect 25688 22720 25740 22772
rect 31392 22720 31444 22772
rect 24952 22584 25004 22636
rect 25136 22627 25188 22636
rect 25136 22593 25145 22627
rect 25145 22593 25179 22627
rect 25179 22593 25188 22627
rect 25136 22584 25188 22593
rect 25504 22584 25556 22636
rect 26240 22627 26292 22636
rect 26240 22593 26249 22627
rect 26249 22593 26283 22627
rect 26283 22593 26292 22627
rect 26240 22584 26292 22593
rect 26424 22584 26476 22636
rect 27988 22652 28040 22704
rect 35072 22652 35124 22704
rect 40776 22652 40828 22704
rect 23940 22559 23992 22568
rect 21272 22448 21324 22500
rect 23940 22525 23949 22559
rect 23949 22525 23983 22559
rect 23983 22525 23992 22559
rect 23940 22516 23992 22525
rect 24216 22448 24268 22500
rect 25596 22516 25648 22568
rect 27344 22516 27396 22568
rect 28632 22584 28684 22636
rect 31852 22584 31904 22636
rect 32680 22584 32732 22636
rect 33508 22584 33560 22636
rect 35900 22584 35952 22636
rect 37740 22627 37792 22636
rect 37740 22593 37749 22627
rect 37749 22593 37783 22627
rect 37783 22593 37792 22627
rect 37740 22584 37792 22593
rect 38384 22627 38436 22636
rect 38384 22593 38393 22627
rect 38393 22593 38427 22627
rect 38427 22593 38436 22627
rect 38384 22584 38436 22593
rect 39764 22584 39816 22636
rect 40960 22627 41012 22636
rect 40960 22593 40969 22627
rect 40969 22593 41003 22627
rect 41003 22593 41012 22627
rect 40960 22584 41012 22593
rect 42524 22584 42576 22636
rect 43352 22584 43404 22636
rect 45652 22652 45704 22704
rect 24952 22448 25004 22500
rect 25780 22448 25832 22500
rect 26240 22448 26292 22500
rect 12440 22380 12492 22389
rect 14464 22380 14516 22432
rect 16028 22423 16080 22432
rect 16028 22389 16037 22423
rect 16037 22389 16071 22423
rect 16071 22389 16080 22423
rect 16028 22380 16080 22389
rect 16580 22380 16632 22432
rect 18512 22380 18564 22432
rect 20628 22380 20680 22432
rect 21180 22423 21232 22432
rect 21180 22389 21189 22423
rect 21189 22389 21223 22423
rect 21223 22389 21232 22423
rect 23204 22423 23256 22432
rect 21180 22380 21232 22389
rect 23204 22389 23213 22423
rect 23213 22389 23247 22423
rect 23247 22389 23256 22423
rect 23204 22380 23256 22389
rect 23756 22380 23808 22432
rect 24032 22380 24084 22432
rect 30104 22559 30156 22568
rect 30104 22525 30113 22559
rect 30113 22525 30147 22559
rect 30147 22525 30156 22559
rect 30104 22516 30156 22525
rect 36544 22516 36596 22568
rect 41880 22559 41932 22568
rect 41880 22525 41889 22559
rect 41889 22525 41923 22559
rect 41923 22525 41932 22559
rect 41880 22516 41932 22525
rect 45284 22559 45336 22568
rect 27804 22380 27856 22432
rect 29092 22380 29144 22432
rect 29644 22380 29696 22432
rect 31576 22423 31628 22432
rect 31576 22389 31585 22423
rect 31585 22389 31619 22423
rect 31619 22389 31628 22423
rect 31576 22380 31628 22389
rect 34060 22423 34112 22432
rect 34060 22389 34069 22423
rect 34069 22389 34103 22423
rect 34103 22389 34112 22423
rect 34060 22380 34112 22389
rect 37740 22380 37792 22432
rect 38752 22380 38804 22432
rect 39212 22423 39264 22432
rect 39212 22389 39221 22423
rect 39221 22389 39255 22423
rect 39255 22389 39264 22423
rect 39212 22380 39264 22389
rect 42524 22423 42576 22432
rect 42524 22389 42533 22423
rect 42533 22389 42567 22423
rect 42567 22389 42576 22423
rect 42524 22380 42576 22389
rect 45284 22525 45293 22559
rect 45293 22525 45327 22559
rect 45327 22525 45336 22559
rect 45284 22516 45336 22525
rect 46572 22448 46624 22500
rect 48320 22695 48372 22704
rect 48320 22661 48329 22695
rect 48329 22661 48363 22695
rect 48363 22661 48372 22695
rect 48320 22652 48372 22661
rect 47676 22516 47728 22568
rect 48596 22559 48648 22568
rect 48596 22525 48605 22559
rect 48605 22525 48639 22559
rect 48639 22525 48648 22559
rect 48596 22516 48648 22525
rect 49148 22516 49200 22568
rect 51908 22584 51960 22636
rect 46848 22380 46900 22432
rect 48044 22448 48096 22500
rect 52276 22448 52328 22500
rect 52000 22423 52052 22432
rect 52000 22389 52009 22423
rect 52009 22389 52043 22423
rect 52043 22389 52052 22423
rect 52000 22380 52052 22389
rect 8174 22278 8226 22330
rect 8238 22278 8290 22330
rect 8302 22278 8354 22330
rect 8366 22278 8418 22330
rect 8430 22278 8482 22330
rect 22622 22278 22674 22330
rect 22686 22278 22738 22330
rect 22750 22278 22802 22330
rect 22814 22278 22866 22330
rect 22878 22278 22930 22330
rect 37070 22278 37122 22330
rect 37134 22278 37186 22330
rect 37198 22278 37250 22330
rect 37262 22278 37314 22330
rect 37326 22278 37378 22330
rect 51518 22278 51570 22330
rect 51582 22278 51634 22330
rect 51646 22278 51698 22330
rect 51710 22278 51762 22330
rect 51774 22278 51826 22330
rect 4712 22219 4764 22228
rect 4712 22185 4721 22219
rect 4721 22185 4755 22219
rect 4755 22185 4764 22219
rect 4712 22176 4764 22185
rect 2228 22040 2280 22092
rect 4620 22040 4672 22092
rect 7380 22040 7432 22092
rect 11336 22176 11388 22228
rect 16212 22176 16264 22228
rect 20628 22176 20680 22228
rect 21824 22176 21876 22228
rect 23204 22176 23256 22228
rect 24584 22219 24636 22228
rect 16672 22108 16724 22160
rect 20352 22108 20404 22160
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 16028 22040 16080 22092
rect 17040 22083 17092 22092
rect 17040 22049 17049 22083
rect 17049 22049 17083 22083
rect 17083 22049 17092 22083
rect 17040 22040 17092 22049
rect 17408 22040 17460 22092
rect 18420 22083 18472 22092
rect 18420 22049 18429 22083
rect 18429 22049 18463 22083
rect 18463 22049 18472 22083
rect 18420 22040 18472 22049
rect 18604 22083 18656 22092
rect 18604 22049 18613 22083
rect 18613 22049 18647 22083
rect 18647 22049 18656 22083
rect 18604 22040 18656 22049
rect 20904 22108 20956 22160
rect 23572 22151 23624 22160
rect 23572 22117 23581 22151
rect 23581 22117 23615 22151
rect 23615 22117 23624 22151
rect 23572 22108 23624 22117
rect 24032 22108 24084 22160
rect 24584 22185 24593 22219
rect 24593 22185 24627 22219
rect 24627 22185 24636 22219
rect 24584 22176 24636 22185
rect 28540 22176 28592 22228
rect 30104 22176 30156 22228
rect 39212 22176 39264 22228
rect 45652 22176 45704 22228
rect 49148 22176 49200 22228
rect 49608 22219 49660 22228
rect 49608 22185 49617 22219
rect 49617 22185 49651 22219
rect 49651 22185 49660 22219
rect 49608 22176 49660 22185
rect 25688 22108 25740 22160
rect 27804 22151 27856 22160
rect 27804 22117 27813 22151
rect 27813 22117 27847 22151
rect 27847 22117 27856 22151
rect 27804 22108 27856 22117
rect 28816 22108 28868 22160
rect 40776 22108 40828 22160
rect 44916 22108 44968 22160
rect 21088 22040 21140 22092
rect 2872 21972 2924 22024
rect 3240 22015 3292 22024
rect 3240 21981 3249 22015
rect 3249 21981 3283 22015
rect 3283 21981 3292 22015
rect 3240 21972 3292 21981
rect 16304 22015 16356 22024
rect 16304 21981 16313 22015
rect 16313 21981 16347 22015
rect 16347 21981 16356 22015
rect 16304 21972 16356 21981
rect 6184 21947 6236 21956
rect 6184 21913 6193 21947
rect 6193 21913 6227 21947
rect 6227 21913 6236 21947
rect 6184 21904 6236 21913
rect 7656 21904 7708 21956
rect 8024 21904 8076 21956
rect 9680 21947 9732 21956
rect 9680 21913 9689 21947
rect 9689 21913 9723 21947
rect 9723 21913 9732 21947
rect 9680 21904 9732 21913
rect 10140 21904 10192 21956
rect 12440 21904 12492 21956
rect 13728 21904 13780 21956
rect 2872 21836 2924 21888
rect 3700 21836 3752 21888
rect 6736 21836 6788 21888
rect 8944 21836 8996 21888
rect 11152 21879 11204 21888
rect 11152 21845 11161 21879
rect 11161 21845 11195 21879
rect 11195 21845 11204 21879
rect 11152 21836 11204 21845
rect 11612 21879 11664 21888
rect 11612 21845 11621 21879
rect 11621 21845 11655 21879
rect 11655 21845 11664 21879
rect 11612 21836 11664 21845
rect 14096 21879 14148 21888
rect 14096 21845 14105 21879
rect 14105 21845 14139 21879
rect 14139 21845 14148 21879
rect 14096 21836 14148 21845
rect 15016 21904 15068 21956
rect 15844 21904 15896 21956
rect 16488 21972 16540 22024
rect 19340 21972 19392 22024
rect 19616 22015 19668 22024
rect 19616 21981 19625 22015
rect 19625 21981 19659 22015
rect 19659 21981 19668 22015
rect 19616 21972 19668 21981
rect 19156 21904 19208 21956
rect 20628 21972 20680 22024
rect 22468 22015 22520 22024
rect 20168 21836 20220 21888
rect 20996 21836 21048 21888
rect 21088 21879 21140 21888
rect 21088 21845 21097 21879
rect 21097 21845 21131 21879
rect 21131 21845 21140 21879
rect 22468 21981 22477 22015
rect 22477 21981 22511 22015
rect 22511 21981 22520 22015
rect 22468 21972 22520 21981
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 25780 22040 25832 22092
rect 24400 21972 24452 22024
rect 24952 21972 25004 22024
rect 25596 22015 25648 22024
rect 25596 21981 25605 22015
rect 25605 21981 25639 22015
rect 25639 21981 25648 22015
rect 25596 21972 25648 21981
rect 26056 22015 26108 22024
rect 26056 21981 26065 22015
rect 26065 21981 26099 22015
rect 26099 21981 26108 22015
rect 26056 21972 26108 21981
rect 21824 21947 21876 21956
rect 21824 21913 21833 21947
rect 21833 21913 21867 21947
rect 21867 21913 21876 21947
rect 21824 21904 21876 21913
rect 23848 21904 23900 21956
rect 24216 21904 24268 21956
rect 25964 21904 26016 21956
rect 26516 21972 26568 22024
rect 29736 22040 29788 22092
rect 31576 22083 31628 22092
rect 31576 22049 31585 22083
rect 31585 22049 31619 22083
rect 31619 22049 31628 22083
rect 31576 22040 31628 22049
rect 33876 22040 33928 22092
rect 27160 21972 27212 22024
rect 21088 21836 21140 21845
rect 24492 21836 24544 21888
rect 24860 21879 24912 21888
rect 24860 21845 24869 21879
rect 24869 21845 24903 21879
rect 24903 21845 24912 21879
rect 24860 21836 24912 21845
rect 25504 21879 25556 21888
rect 25504 21845 25513 21879
rect 25513 21845 25547 21879
rect 25547 21845 25556 21879
rect 25504 21836 25556 21845
rect 26148 21879 26200 21888
rect 26148 21845 26157 21879
rect 26157 21845 26191 21879
rect 26191 21845 26200 21879
rect 26148 21836 26200 21845
rect 27344 21836 27396 21888
rect 27988 22015 28040 22024
rect 27988 21981 27997 22015
rect 27997 21981 28031 22015
rect 28031 21981 28040 22015
rect 27988 21972 28040 21981
rect 28264 21972 28316 22024
rect 29000 22015 29052 22024
rect 29000 21981 29009 22015
rect 29009 21981 29043 22015
rect 29043 21981 29052 22015
rect 29000 21972 29052 21981
rect 30472 22015 30524 22024
rect 28356 21904 28408 21956
rect 30472 21981 30481 22015
rect 30481 21981 30515 22015
rect 30515 21981 30524 22015
rect 30472 21972 30524 21981
rect 34152 22015 34204 22024
rect 31300 21904 31352 21956
rect 34152 21981 34161 22015
rect 34161 21981 34195 22015
rect 34195 21981 34204 22015
rect 34152 21972 34204 21981
rect 35900 21972 35952 22024
rect 36728 22015 36780 22024
rect 36728 21981 36737 22015
rect 36737 21981 36771 22015
rect 36771 21981 36780 22015
rect 36728 21972 36780 21981
rect 39304 21972 39356 22024
rect 40040 22015 40092 22024
rect 40040 21981 40049 22015
rect 40049 21981 40083 22015
rect 40083 21981 40092 22015
rect 40040 21972 40092 21981
rect 43444 21972 43496 22024
rect 37740 21904 37792 21956
rect 29460 21836 29512 21888
rect 30564 21879 30616 21888
rect 30564 21845 30573 21879
rect 30573 21845 30607 21879
rect 30607 21845 30616 21879
rect 30564 21836 30616 21845
rect 32312 21879 32364 21888
rect 32312 21845 32321 21879
rect 32321 21845 32355 21879
rect 32355 21845 32364 21879
rect 32312 21836 32364 21845
rect 36912 21836 36964 21888
rect 38568 21836 38620 21888
rect 39488 21836 39540 21888
rect 45284 22040 45336 22092
rect 47216 22040 47268 22092
rect 48320 22083 48372 22092
rect 48320 22049 48329 22083
rect 48329 22049 48363 22083
rect 48363 22049 48372 22083
rect 48320 22040 48372 22049
rect 44088 21972 44140 22024
rect 45376 22015 45428 22024
rect 45376 21981 45385 22015
rect 45385 21981 45419 22015
rect 45419 21981 45428 22015
rect 45376 21972 45428 21981
rect 46204 21972 46256 22024
rect 47768 21972 47820 22024
rect 50160 21972 50212 22024
rect 50620 22040 50672 22092
rect 50712 21972 50764 22024
rect 45284 21904 45336 21956
rect 48412 21904 48464 21956
rect 55128 21972 55180 22024
rect 51908 21904 51960 21956
rect 44180 21836 44232 21888
rect 45008 21879 45060 21888
rect 45008 21845 45017 21879
rect 45017 21845 45051 21879
rect 45051 21845 45060 21879
rect 45008 21836 45060 21845
rect 45744 21836 45796 21888
rect 46572 21879 46624 21888
rect 46572 21845 46581 21879
rect 46581 21845 46615 21879
rect 46615 21845 46624 21879
rect 46572 21836 46624 21845
rect 47584 21879 47636 21888
rect 47584 21845 47593 21879
rect 47593 21845 47627 21879
rect 47627 21845 47636 21879
rect 47584 21836 47636 21845
rect 48596 21879 48648 21888
rect 48596 21845 48605 21879
rect 48605 21845 48639 21879
rect 48639 21845 48648 21879
rect 48596 21836 48648 21845
rect 49240 21879 49292 21888
rect 49240 21845 49249 21879
rect 49249 21845 49283 21879
rect 49283 21845 49292 21879
rect 49240 21836 49292 21845
rect 49976 21836 50028 21888
rect 52368 21836 52420 21888
rect 55588 21879 55640 21888
rect 55588 21845 55597 21879
rect 55597 21845 55631 21879
rect 55631 21845 55640 21879
rect 55588 21836 55640 21845
rect 15398 21734 15450 21786
rect 15462 21734 15514 21786
rect 15526 21734 15578 21786
rect 15590 21734 15642 21786
rect 15654 21734 15706 21786
rect 29846 21734 29898 21786
rect 29910 21734 29962 21786
rect 29974 21734 30026 21786
rect 30038 21734 30090 21786
rect 30102 21734 30154 21786
rect 44294 21734 44346 21786
rect 44358 21734 44410 21786
rect 44422 21734 44474 21786
rect 44486 21734 44538 21786
rect 44550 21734 44602 21786
rect 3976 21632 4028 21684
rect 2872 21564 2924 21616
rect 5448 21564 5500 21616
rect 5908 21564 5960 21616
rect 6184 21632 6236 21684
rect 11796 21675 11848 21684
rect 6736 21564 6788 21616
rect 7104 21564 7156 21616
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 13176 21632 13228 21684
rect 17960 21632 18012 21684
rect 20168 21632 20220 21684
rect 21088 21632 21140 21684
rect 9404 21564 9456 21616
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 10416 21539 10468 21548
rect 5816 21496 5868 21505
rect 10416 21505 10425 21539
rect 10425 21505 10459 21539
rect 10459 21505 10468 21539
rect 10416 21496 10468 21505
rect 3332 21471 3384 21480
rect 3332 21437 3341 21471
rect 3341 21437 3375 21471
rect 3375 21437 3384 21471
rect 3332 21428 3384 21437
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 4344 21428 4396 21480
rect 5080 21292 5132 21344
rect 6736 21428 6788 21480
rect 16304 21564 16356 21616
rect 17132 21607 17184 21616
rect 17132 21573 17141 21607
rect 17141 21573 17175 21607
rect 17175 21573 17184 21607
rect 17132 21564 17184 21573
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 11796 21496 11848 21548
rect 15016 21496 15068 21548
rect 15752 21539 15804 21548
rect 15752 21505 15761 21539
rect 15761 21505 15795 21539
rect 15795 21505 15804 21539
rect 15752 21496 15804 21505
rect 16396 21496 16448 21548
rect 18696 21539 18748 21548
rect 18696 21505 18705 21539
rect 18705 21505 18739 21539
rect 18739 21505 18748 21539
rect 18696 21496 18748 21505
rect 19616 21564 19668 21616
rect 24952 21632 25004 21684
rect 25596 21632 25648 21684
rect 27804 21632 27856 21684
rect 27896 21632 27948 21684
rect 25504 21564 25556 21616
rect 26056 21564 26108 21616
rect 26884 21564 26936 21616
rect 27528 21564 27580 21616
rect 27620 21564 27672 21616
rect 30196 21607 30248 21616
rect 30196 21573 30205 21607
rect 30205 21573 30239 21607
rect 30239 21573 30248 21607
rect 30196 21564 30248 21573
rect 22284 21539 22336 21548
rect 15292 21428 15344 21480
rect 18328 21428 18380 21480
rect 10968 21360 11020 21412
rect 17776 21360 17828 21412
rect 19248 21428 19300 21480
rect 19800 21471 19852 21480
rect 19156 21360 19208 21412
rect 19800 21437 19809 21471
rect 19809 21437 19843 21471
rect 19843 21437 19852 21471
rect 19800 21428 19852 21437
rect 20720 21428 20772 21480
rect 7196 21292 7248 21344
rect 12992 21292 13044 21344
rect 15752 21292 15804 21344
rect 17408 21335 17460 21344
rect 17408 21301 17417 21335
rect 17417 21301 17451 21335
rect 17451 21301 17460 21335
rect 17408 21292 17460 21301
rect 20352 21360 20404 21412
rect 22284 21505 22293 21539
rect 22293 21505 22327 21539
rect 22327 21505 22336 21539
rect 22284 21496 22336 21505
rect 23296 21539 23348 21548
rect 23296 21505 23305 21539
rect 23305 21505 23339 21539
rect 23339 21505 23348 21539
rect 23296 21496 23348 21505
rect 24860 21496 24912 21548
rect 26240 21539 26292 21548
rect 26240 21505 26249 21539
rect 26249 21505 26283 21539
rect 26283 21505 26292 21539
rect 26240 21496 26292 21505
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 27252 21496 27304 21548
rect 27896 21496 27948 21548
rect 28172 21539 28224 21548
rect 28172 21505 28181 21539
rect 28181 21505 28215 21539
rect 28215 21505 28224 21539
rect 28172 21496 28224 21505
rect 31576 21496 31628 21548
rect 32864 21539 32916 21548
rect 32864 21505 32873 21539
rect 32873 21505 32907 21539
rect 32907 21505 32916 21539
rect 32864 21496 32916 21505
rect 35440 21632 35492 21684
rect 36268 21675 36320 21684
rect 36268 21641 36277 21675
rect 36277 21641 36311 21675
rect 36311 21641 36320 21675
rect 36268 21632 36320 21641
rect 39764 21675 39816 21684
rect 39764 21641 39773 21675
rect 39773 21641 39807 21675
rect 39807 21641 39816 21675
rect 39764 21632 39816 21641
rect 23664 21428 23716 21480
rect 24952 21428 25004 21480
rect 25872 21360 25924 21412
rect 27068 21428 27120 21480
rect 26516 21360 26568 21412
rect 26884 21360 26936 21412
rect 28080 21428 28132 21480
rect 30472 21428 30524 21480
rect 34520 21496 34572 21548
rect 35624 21496 35676 21548
rect 37004 21496 37056 21548
rect 38568 21564 38620 21616
rect 38016 21539 38068 21548
rect 38016 21505 38025 21539
rect 38025 21505 38059 21539
rect 38059 21505 38068 21539
rect 38016 21496 38068 21505
rect 40408 21539 40460 21548
rect 40408 21505 40417 21539
rect 40417 21505 40451 21539
rect 40451 21505 40460 21539
rect 40408 21496 40460 21505
rect 45376 21632 45428 21684
rect 47492 21632 47544 21684
rect 45652 21564 45704 21616
rect 49516 21632 49568 21684
rect 49608 21632 49660 21684
rect 48596 21564 48648 21616
rect 49148 21564 49200 21616
rect 45008 21496 45060 21548
rect 47676 21496 47728 21548
rect 47768 21496 47820 21548
rect 48412 21539 48464 21548
rect 36820 21428 36872 21480
rect 39304 21428 39356 21480
rect 42616 21471 42668 21480
rect 42616 21437 42625 21471
rect 42625 21437 42659 21471
rect 42659 21437 42668 21471
rect 42616 21428 42668 21437
rect 42708 21428 42760 21480
rect 27344 21403 27396 21412
rect 27344 21369 27353 21403
rect 27353 21369 27387 21403
rect 27387 21369 27396 21403
rect 27344 21360 27396 21369
rect 27528 21360 27580 21412
rect 29368 21360 29420 21412
rect 21272 21292 21324 21344
rect 21640 21292 21692 21344
rect 22468 21292 22520 21344
rect 24952 21292 25004 21344
rect 26240 21292 26292 21344
rect 27620 21292 27672 21344
rect 27804 21292 27856 21344
rect 28816 21292 28868 21344
rect 31852 21360 31904 21412
rect 43628 21360 43680 21412
rect 29828 21292 29880 21344
rect 32036 21292 32088 21344
rect 33416 21335 33468 21344
rect 33416 21301 33425 21335
rect 33425 21301 33459 21335
rect 33459 21301 33468 21335
rect 33416 21292 33468 21301
rect 35808 21292 35860 21344
rect 43444 21292 43496 21344
rect 47400 21428 47452 21480
rect 47768 21360 47820 21412
rect 47400 21292 47452 21344
rect 48412 21505 48421 21539
rect 48421 21505 48455 21539
rect 48455 21505 48464 21539
rect 48412 21496 48464 21505
rect 50712 21496 50764 21548
rect 53104 21496 53156 21548
rect 56692 21496 56744 21548
rect 49332 21428 49384 21480
rect 52000 21428 52052 21480
rect 54300 21428 54352 21480
rect 55128 21428 55180 21480
rect 55772 21428 55824 21480
rect 49056 21292 49108 21344
rect 52828 21335 52880 21344
rect 52828 21301 52837 21335
rect 52837 21301 52871 21335
rect 52871 21301 52880 21335
rect 52828 21292 52880 21301
rect 55496 21292 55548 21344
rect 8174 21190 8226 21242
rect 8238 21190 8290 21242
rect 8302 21190 8354 21242
rect 8366 21190 8418 21242
rect 8430 21190 8482 21242
rect 22622 21190 22674 21242
rect 22686 21190 22738 21242
rect 22750 21190 22802 21242
rect 22814 21190 22866 21242
rect 22878 21190 22930 21242
rect 37070 21190 37122 21242
rect 37134 21190 37186 21242
rect 37198 21190 37250 21242
rect 37262 21190 37314 21242
rect 37326 21190 37378 21242
rect 51518 21190 51570 21242
rect 51582 21190 51634 21242
rect 51646 21190 51698 21242
rect 51710 21190 51762 21242
rect 51774 21190 51826 21242
rect 2964 21088 3016 21140
rect 3608 21088 3660 21140
rect 6736 21088 6788 21140
rect 7012 21088 7064 21140
rect 5448 21020 5500 21072
rect 7656 21020 7708 21072
rect 3240 20952 3292 21004
rect 3976 20952 4028 21004
rect 6552 20952 6604 21004
rect 10324 20952 10376 21004
rect 16120 21088 16172 21140
rect 19432 21131 19484 21140
rect 19432 21097 19441 21131
rect 19441 21097 19475 21131
rect 19475 21097 19484 21131
rect 19432 21088 19484 21097
rect 20536 21131 20588 21140
rect 20536 21097 20545 21131
rect 20545 21097 20579 21131
rect 20579 21097 20588 21131
rect 20536 21088 20588 21097
rect 22100 21131 22152 21140
rect 22100 21097 22109 21131
rect 22109 21097 22143 21131
rect 22143 21097 22152 21131
rect 22100 21088 22152 21097
rect 23664 21131 23716 21140
rect 23664 21097 23673 21131
rect 23673 21097 23707 21131
rect 23707 21097 23716 21131
rect 23664 21088 23716 21097
rect 24400 21131 24452 21140
rect 24400 21097 24409 21131
rect 24409 21097 24443 21131
rect 24443 21097 24452 21131
rect 24400 21088 24452 21097
rect 24952 21088 25004 21140
rect 27068 21088 27120 21140
rect 27252 21131 27304 21140
rect 27252 21097 27261 21131
rect 27261 21097 27295 21131
rect 27295 21097 27304 21131
rect 27252 21088 27304 21097
rect 27988 21088 28040 21140
rect 31300 21131 31352 21140
rect 31300 21097 31309 21131
rect 31309 21097 31343 21131
rect 31343 21097 31352 21131
rect 31300 21088 31352 21097
rect 33508 21131 33560 21140
rect 33508 21097 33517 21131
rect 33517 21097 33551 21131
rect 33551 21097 33560 21131
rect 33508 21088 33560 21097
rect 36360 21131 36412 21140
rect 36360 21097 36369 21131
rect 36369 21097 36403 21131
rect 36403 21097 36412 21131
rect 36360 21088 36412 21097
rect 37832 21131 37884 21140
rect 37832 21097 37841 21131
rect 37841 21097 37875 21131
rect 37875 21097 37884 21131
rect 37832 21088 37884 21097
rect 42984 21088 43036 21140
rect 46204 21088 46256 21140
rect 47216 21131 47268 21140
rect 47216 21097 47225 21131
rect 47225 21097 47259 21131
rect 47259 21097 47268 21131
rect 47216 21088 47268 21097
rect 47492 21088 47544 21140
rect 49332 21131 49384 21140
rect 49332 21097 49341 21131
rect 49341 21097 49375 21131
rect 49375 21097 49384 21131
rect 49332 21088 49384 21097
rect 50620 21131 50672 21140
rect 50620 21097 50629 21131
rect 50629 21097 50663 21131
rect 50663 21097 50672 21131
rect 50620 21088 50672 21097
rect 17132 21020 17184 21072
rect 19616 21020 19668 21072
rect 12532 20952 12584 21004
rect 4988 20884 5040 20936
rect 9404 20927 9456 20936
rect 9404 20893 9413 20927
rect 9413 20893 9447 20927
rect 9447 20893 9456 20927
rect 9404 20884 9456 20893
rect 13544 20884 13596 20936
rect 17040 20952 17092 21004
rect 20260 20952 20312 21004
rect 15200 20884 15252 20936
rect 16488 20884 16540 20936
rect 18696 20884 18748 20936
rect 20352 20927 20404 20936
rect 20352 20893 20361 20927
rect 20361 20893 20395 20927
rect 20395 20893 20404 20927
rect 20352 20884 20404 20893
rect 21088 21020 21140 21072
rect 21548 21063 21600 21072
rect 21272 20995 21324 21004
rect 21272 20961 21281 20995
rect 21281 20961 21315 20995
rect 21315 20961 21324 20995
rect 21272 20952 21324 20961
rect 21548 21029 21557 21063
rect 21557 21029 21591 21063
rect 21591 21029 21600 21063
rect 21548 21020 21600 21029
rect 21824 21020 21876 21072
rect 23848 21020 23900 21072
rect 22192 20884 22244 20936
rect 22284 20884 22336 20936
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 23848 20884 23900 20893
rect 4252 20748 4304 20800
rect 10784 20748 10836 20800
rect 14648 20816 14700 20868
rect 26148 21020 26200 21072
rect 26516 21063 26568 21072
rect 25228 20884 25280 20936
rect 26240 20884 26292 20936
rect 26516 21029 26525 21063
rect 26525 21029 26559 21063
rect 26559 21029 26568 21063
rect 26516 21020 26568 21029
rect 27896 21020 27948 21072
rect 27344 20952 27396 21004
rect 29000 21020 29052 21072
rect 29276 20952 29328 21004
rect 29828 20995 29880 21004
rect 29828 20961 29837 20995
rect 29837 20961 29871 20995
rect 29871 20961 29880 20995
rect 29828 20952 29880 20961
rect 31760 20995 31812 21004
rect 31760 20961 31769 20995
rect 31769 20961 31803 20995
rect 31803 20961 31812 20995
rect 32036 20995 32088 21004
rect 31760 20952 31812 20961
rect 32036 20961 32045 20995
rect 32045 20961 32079 20995
rect 32079 20961 32088 20995
rect 32036 20952 32088 20961
rect 32404 20952 32456 21004
rect 27436 20927 27488 20936
rect 27436 20893 27445 20927
rect 27445 20893 27479 20927
rect 27479 20893 27488 20927
rect 27436 20884 27488 20893
rect 28724 20884 28776 20936
rect 34612 20884 34664 20936
rect 35532 21020 35584 21072
rect 40592 21020 40644 21072
rect 42616 21020 42668 21072
rect 42708 20952 42760 21004
rect 43996 21020 44048 21072
rect 44272 21020 44324 21072
rect 44824 21020 44876 21072
rect 43628 20995 43680 21004
rect 43628 20961 43637 20995
rect 43637 20961 43671 20995
rect 43671 20961 43680 20995
rect 43628 20952 43680 20961
rect 46848 21020 46900 21072
rect 36544 20927 36596 20936
rect 15200 20791 15252 20800
rect 15200 20757 15209 20791
rect 15209 20757 15243 20791
rect 15243 20757 15252 20791
rect 15200 20748 15252 20757
rect 16488 20748 16540 20800
rect 18420 20791 18472 20800
rect 18420 20757 18429 20791
rect 18429 20757 18463 20791
rect 18463 20757 18472 20791
rect 18420 20748 18472 20757
rect 20444 20748 20496 20800
rect 29736 20816 29788 20868
rect 30564 20816 30616 20868
rect 33416 20816 33468 20868
rect 25688 20791 25740 20800
rect 25688 20757 25697 20791
rect 25697 20757 25731 20791
rect 25731 20757 25740 20791
rect 25688 20748 25740 20757
rect 29092 20748 29144 20800
rect 32864 20748 32916 20800
rect 36544 20893 36553 20927
rect 36553 20893 36587 20927
rect 36587 20893 36596 20927
rect 36544 20884 36596 20893
rect 37004 20927 37056 20936
rect 37004 20893 37013 20927
rect 37013 20893 37047 20927
rect 37047 20893 37056 20927
rect 37004 20884 37056 20893
rect 37924 20884 37976 20936
rect 39948 20927 40000 20936
rect 39948 20893 39957 20927
rect 39957 20893 39991 20927
rect 39991 20893 40000 20927
rect 39948 20884 40000 20893
rect 40040 20884 40092 20936
rect 44180 20884 44232 20936
rect 36544 20748 36596 20800
rect 37924 20748 37976 20800
rect 38476 20748 38528 20800
rect 41328 20748 41380 20800
rect 42432 20816 42484 20868
rect 44088 20816 44140 20868
rect 44732 20816 44784 20868
rect 44916 20816 44968 20868
rect 45744 20884 45796 20936
rect 47400 20927 47452 20936
rect 47400 20893 47409 20927
rect 47409 20893 47443 20927
rect 47443 20893 47452 20927
rect 47400 20884 47452 20893
rect 47676 20927 47728 20936
rect 47676 20893 47685 20927
rect 47685 20893 47719 20927
rect 47719 20893 47728 20927
rect 47676 20884 47728 20893
rect 47768 20927 47820 20936
rect 47768 20893 47777 20927
rect 47777 20893 47811 20927
rect 47811 20893 47820 20927
rect 48412 20927 48464 20936
rect 47768 20884 47820 20893
rect 48412 20893 48421 20927
rect 48421 20893 48455 20927
rect 48455 20893 48464 20927
rect 48412 20884 48464 20893
rect 49240 20952 49292 21004
rect 50344 21020 50396 21072
rect 44272 20748 44324 20800
rect 44640 20748 44692 20800
rect 46480 20748 46532 20800
rect 49056 20816 49108 20868
rect 50160 20927 50212 20936
rect 50160 20893 50169 20927
rect 50169 20893 50203 20927
rect 50203 20893 50212 20927
rect 50160 20884 50212 20893
rect 50436 20927 50488 20936
rect 50436 20893 50445 20927
rect 50445 20893 50479 20927
rect 50479 20893 50488 20927
rect 50436 20884 50488 20893
rect 55496 21088 55548 21140
rect 55772 21131 55824 21140
rect 55772 21097 55781 21131
rect 55781 21097 55815 21131
rect 55815 21097 55824 21131
rect 55772 21088 55824 21097
rect 52000 20952 52052 21004
rect 52368 20952 52420 21004
rect 49516 20859 49568 20868
rect 49516 20825 49525 20859
rect 49525 20825 49559 20859
rect 49559 20825 49568 20859
rect 49516 20816 49568 20825
rect 50068 20816 50120 20868
rect 51264 20927 51316 20936
rect 51264 20893 51273 20927
rect 51273 20893 51307 20927
rect 51307 20893 51316 20927
rect 51264 20884 51316 20893
rect 52000 20859 52052 20868
rect 48872 20748 48924 20800
rect 52000 20825 52009 20859
rect 52009 20825 52043 20859
rect 52043 20825 52052 20859
rect 52000 20816 52052 20825
rect 53656 20952 53708 21004
rect 53288 20884 53340 20936
rect 54116 20927 54168 20936
rect 54116 20893 54125 20927
rect 54125 20893 54159 20927
rect 54159 20893 54168 20927
rect 55496 20927 55548 20936
rect 54116 20884 54168 20893
rect 55496 20893 55505 20927
rect 55505 20893 55539 20927
rect 55539 20893 55548 20927
rect 55496 20884 55548 20893
rect 56692 20927 56744 20936
rect 56692 20893 56701 20927
rect 56701 20893 56735 20927
rect 56735 20893 56744 20927
rect 56692 20884 56744 20893
rect 57336 20816 57388 20868
rect 53288 20748 53340 20800
rect 53472 20791 53524 20800
rect 53472 20757 53481 20791
rect 53481 20757 53515 20791
rect 53515 20757 53524 20791
rect 53472 20748 53524 20757
rect 15398 20646 15450 20698
rect 15462 20646 15514 20698
rect 15526 20646 15578 20698
rect 15590 20646 15642 20698
rect 15654 20646 15706 20698
rect 29846 20646 29898 20698
rect 29910 20646 29962 20698
rect 29974 20646 30026 20698
rect 30038 20646 30090 20698
rect 30102 20646 30154 20698
rect 44294 20646 44346 20698
rect 44358 20646 44410 20698
rect 44422 20646 44474 20698
rect 44486 20646 44538 20698
rect 44550 20646 44602 20698
rect 2964 20587 3016 20596
rect 2964 20553 2973 20587
rect 2973 20553 3007 20587
rect 3007 20553 3016 20587
rect 2964 20544 3016 20553
rect 3608 20587 3660 20596
rect 3608 20553 3617 20587
rect 3617 20553 3651 20587
rect 3651 20553 3660 20587
rect 3608 20544 3660 20553
rect 4804 20544 4856 20596
rect 7104 20544 7156 20596
rect 7380 20544 7432 20596
rect 9128 20587 9180 20596
rect 9128 20553 9137 20587
rect 9137 20553 9171 20587
rect 9171 20553 9180 20587
rect 9128 20544 9180 20553
rect 11796 20544 11848 20596
rect 14464 20587 14516 20596
rect 14464 20553 14473 20587
rect 14473 20553 14507 20587
rect 14507 20553 14516 20587
rect 14464 20544 14516 20553
rect 15200 20544 15252 20596
rect 19340 20544 19392 20596
rect 20904 20544 20956 20596
rect 21364 20544 21416 20596
rect 24124 20544 24176 20596
rect 7840 20519 7892 20528
rect 7840 20485 7849 20519
rect 7849 20485 7883 20519
rect 7883 20485 7892 20519
rect 7840 20476 7892 20485
rect 9772 20476 9824 20528
rect 16764 20476 16816 20528
rect 2136 20408 2188 20460
rect 2780 20451 2832 20460
rect 2780 20417 2789 20451
rect 2789 20417 2823 20451
rect 2823 20417 2832 20451
rect 2780 20408 2832 20417
rect 6368 20408 6420 20460
rect 7012 20408 7064 20460
rect 7656 20408 7708 20460
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 11428 20408 11480 20460
rect 14004 20451 14056 20460
rect 14004 20417 14013 20451
rect 14013 20417 14047 20451
rect 14047 20417 14056 20451
rect 14004 20408 14056 20417
rect 16396 20408 16448 20460
rect 16488 20408 16540 20460
rect 17868 20476 17920 20528
rect 23020 20476 23072 20528
rect 25688 20519 25740 20528
rect 25688 20485 25697 20519
rect 25697 20485 25731 20519
rect 25731 20485 25740 20519
rect 25688 20476 25740 20485
rect 26148 20544 26200 20596
rect 28356 20544 28408 20596
rect 27896 20476 27948 20528
rect 28264 20476 28316 20528
rect 22192 20451 22244 20460
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 25964 20451 26016 20460
rect 25964 20417 25973 20451
rect 25973 20417 26007 20451
rect 26007 20417 26016 20451
rect 27620 20451 27672 20460
rect 25964 20408 26016 20417
rect 27620 20417 27629 20451
rect 27629 20417 27663 20451
rect 27663 20417 27672 20451
rect 27620 20408 27672 20417
rect 28080 20408 28132 20460
rect 29460 20544 29512 20596
rect 30104 20476 30156 20528
rect 32404 20519 32456 20528
rect 32404 20485 32413 20519
rect 32413 20485 32447 20519
rect 32447 20485 32456 20519
rect 32404 20476 32456 20485
rect 32956 20476 33008 20528
rect 35808 20476 35860 20528
rect 34520 20451 34572 20460
rect 34520 20417 34529 20451
rect 34529 20417 34563 20451
rect 34563 20417 34572 20451
rect 34520 20408 34572 20417
rect 39948 20544 40000 20596
rect 38752 20476 38804 20528
rect 37464 20408 37516 20460
rect 40316 20451 40368 20460
rect 40316 20417 40325 20451
rect 40325 20417 40359 20451
rect 40359 20417 40368 20451
rect 40316 20408 40368 20417
rect 40592 20408 40644 20460
rect 43352 20476 43404 20528
rect 42984 20408 43036 20460
rect 43996 20451 44048 20460
rect 43996 20417 44005 20451
rect 44005 20417 44039 20451
rect 44039 20417 44048 20451
rect 43996 20408 44048 20417
rect 44640 20451 44692 20460
rect 44640 20417 44649 20451
rect 44649 20417 44683 20451
rect 44683 20417 44692 20451
rect 44640 20408 44692 20417
rect 45744 20408 45796 20460
rect 46296 20451 46348 20460
rect 46296 20417 46305 20451
rect 46305 20417 46339 20451
rect 46339 20417 46348 20451
rect 46296 20408 46348 20417
rect 47492 20408 47544 20460
rect 47768 20408 47820 20460
rect 49976 20544 50028 20596
rect 50344 20544 50396 20596
rect 49608 20476 49660 20528
rect 52000 20544 52052 20596
rect 52828 20544 52880 20596
rect 53288 20587 53340 20596
rect 53288 20553 53297 20587
rect 53297 20553 53331 20587
rect 53331 20553 53340 20587
rect 53288 20544 53340 20553
rect 54116 20544 54168 20596
rect 53472 20476 53524 20528
rect 52460 20408 52512 20460
rect 2872 20340 2924 20392
rect 3792 20340 3844 20392
rect 11796 20383 11848 20392
rect 11796 20349 11805 20383
rect 11805 20349 11839 20383
rect 11839 20349 11848 20383
rect 11796 20340 11848 20349
rect 7288 20272 7340 20324
rect 8760 20204 8812 20256
rect 13544 20272 13596 20324
rect 17040 20340 17092 20392
rect 18328 20340 18380 20392
rect 21272 20340 21324 20392
rect 31024 20340 31076 20392
rect 19156 20272 19208 20324
rect 39488 20340 39540 20392
rect 43628 20340 43680 20392
rect 45376 20383 45428 20392
rect 45376 20349 45385 20383
rect 45385 20349 45419 20383
rect 45419 20349 45428 20383
rect 45376 20340 45428 20349
rect 49700 20340 49752 20392
rect 50528 20340 50580 20392
rect 51356 20383 51408 20392
rect 51356 20349 51365 20383
rect 51365 20349 51399 20383
rect 51399 20349 51408 20383
rect 51356 20340 51408 20349
rect 53748 20340 53800 20392
rect 13176 20204 13228 20256
rect 15568 20247 15620 20256
rect 15568 20213 15577 20247
rect 15577 20213 15611 20247
rect 15611 20213 15620 20247
rect 15568 20204 15620 20213
rect 16764 20247 16816 20256
rect 16764 20213 16773 20247
rect 16773 20213 16807 20247
rect 16807 20213 16816 20247
rect 16764 20204 16816 20213
rect 17776 20247 17828 20256
rect 17776 20213 17785 20247
rect 17785 20213 17819 20247
rect 17819 20213 17828 20247
rect 17776 20204 17828 20213
rect 21272 20204 21324 20256
rect 23296 20204 23348 20256
rect 23848 20204 23900 20256
rect 25688 20204 25740 20256
rect 27436 20204 27488 20256
rect 34336 20204 34388 20256
rect 34612 20204 34664 20256
rect 35072 20204 35124 20256
rect 39396 20204 39448 20256
rect 40132 20204 40184 20256
rect 41236 20247 41288 20256
rect 41236 20213 41245 20247
rect 41245 20213 41279 20247
rect 41279 20213 41288 20247
rect 41236 20204 41288 20213
rect 41788 20247 41840 20256
rect 41788 20213 41797 20247
rect 41797 20213 41831 20247
rect 41831 20213 41840 20247
rect 41788 20204 41840 20213
rect 42432 20204 42484 20256
rect 43076 20204 43128 20256
rect 48412 20272 48464 20324
rect 44732 20204 44784 20256
rect 46572 20204 46624 20256
rect 48688 20247 48740 20256
rect 48688 20213 48697 20247
rect 48697 20213 48731 20247
rect 48731 20213 48740 20247
rect 48688 20204 48740 20213
rect 52092 20272 52144 20324
rect 53840 20272 53892 20324
rect 50436 20204 50488 20256
rect 52920 20204 52972 20256
rect 55220 20204 55272 20256
rect 8174 20102 8226 20154
rect 8238 20102 8290 20154
rect 8302 20102 8354 20154
rect 8366 20102 8418 20154
rect 8430 20102 8482 20154
rect 22622 20102 22674 20154
rect 22686 20102 22738 20154
rect 22750 20102 22802 20154
rect 22814 20102 22866 20154
rect 22878 20102 22930 20154
rect 37070 20102 37122 20154
rect 37134 20102 37186 20154
rect 37198 20102 37250 20154
rect 37262 20102 37314 20154
rect 37326 20102 37378 20154
rect 51518 20102 51570 20154
rect 51582 20102 51634 20154
rect 51646 20102 51698 20154
rect 51710 20102 51762 20154
rect 51774 20102 51826 20154
rect 7932 20000 7984 20052
rect 10416 20000 10468 20052
rect 13912 20000 13964 20052
rect 17868 20000 17920 20052
rect 20904 20000 20956 20052
rect 3884 19932 3936 19984
rect 5724 19932 5776 19984
rect 2228 19907 2280 19916
rect 2228 19873 2237 19907
rect 2237 19873 2271 19907
rect 2271 19873 2280 19907
rect 2228 19864 2280 19873
rect 2136 19839 2188 19848
rect 2136 19805 2145 19839
rect 2145 19805 2179 19839
rect 2179 19805 2188 19839
rect 2136 19796 2188 19805
rect 3700 19796 3752 19848
rect 9128 19864 9180 19916
rect 11244 19907 11296 19916
rect 11244 19873 11253 19907
rect 11253 19873 11287 19907
rect 11287 19873 11296 19907
rect 11244 19864 11296 19873
rect 15568 19932 15620 19984
rect 18328 19932 18380 19984
rect 22192 19975 22244 19984
rect 22192 19941 22201 19975
rect 22201 19941 22235 19975
rect 22235 19941 22244 19975
rect 22192 19932 22244 19941
rect 22376 20000 22428 20052
rect 25044 20000 25096 20052
rect 25136 20000 25188 20052
rect 30104 20000 30156 20052
rect 32956 20043 33008 20052
rect 32956 20009 32965 20043
rect 32965 20009 32999 20043
rect 32999 20009 33008 20043
rect 32956 20000 33008 20009
rect 12716 19864 12768 19916
rect 16488 19907 16540 19916
rect 6276 19728 6328 19780
rect 7656 19728 7708 19780
rect 9864 19796 9916 19848
rect 10232 19796 10284 19848
rect 10784 19796 10836 19848
rect 14096 19796 14148 19848
rect 16488 19873 16497 19907
rect 16497 19873 16531 19907
rect 16531 19873 16540 19907
rect 16488 19864 16540 19873
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 20444 19864 20496 19916
rect 24860 19864 24912 19916
rect 17132 19839 17184 19848
rect 5632 19660 5684 19712
rect 6368 19660 6420 19712
rect 9772 19660 9824 19712
rect 11060 19728 11112 19780
rect 12532 19728 12584 19780
rect 17132 19805 17141 19839
rect 17141 19805 17175 19839
rect 17175 19805 17184 19839
rect 17132 19796 17184 19805
rect 11612 19660 11664 19712
rect 13360 19660 13412 19712
rect 13544 19703 13596 19712
rect 13544 19669 13553 19703
rect 13553 19669 13587 19703
rect 13587 19669 13596 19703
rect 13544 19660 13596 19669
rect 14372 19660 14424 19712
rect 14556 19703 14608 19712
rect 14556 19669 14565 19703
rect 14565 19669 14599 19703
rect 14599 19669 14608 19703
rect 14556 19660 14608 19669
rect 14740 19660 14792 19712
rect 17408 19728 17460 19780
rect 19616 19796 19668 19848
rect 20904 19796 20956 19848
rect 21272 19839 21324 19848
rect 21272 19805 21281 19839
rect 21281 19805 21315 19839
rect 21315 19805 21324 19839
rect 21272 19796 21324 19805
rect 22468 19796 22520 19848
rect 27620 19932 27672 19984
rect 27896 19932 27948 19984
rect 25688 19864 25740 19916
rect 20628 19728 20680 19780
rect 22284 19728 22336 19780
rect 23020 19728 23072 19780
rect 25872 19796 25924 19848
rect 26240 19796 26292 19848
rect 27896 19796 27948 19848
rect 28264 19796 28316 19848
rect 28816 19839 28868 19848
rect 28816 19805 28825 19839
rect 28825 19805 28859 19839
rect 28859 19805 28868 19839
rect 28816 19796 28868 19805
rect 30472 19796 30524 19848
rect 30656 19839 30708 19848
rect 30656 19805 30665 19839
rect 30665 19805 30699 19839
rect 30699 19805 30708 19839
rect 30656 19796 30708 19805
rect 25136 19728 25188 19780
rect 27804 19771 27856 19780
rect 19248 19660 19300 19712
rect 19892 19703 19944 19712
rect 19892 19669 19901 19703
rect 19901 19669 19935 19703
rect 19935 19669 19944 19703
rect 19892 19660 19944 19669
rect 23756 19703 23808 19712
rect 23756 19669 23765 19703
rect 23765 19669 23799 19703
rect 23799 19669 23808 19703
rect 23756 19660 23808 19669
rect 27344 19703 27396 19712
rect 27344 19669 27353 19703
rect 27353 19669 27387 19703
rect 27387 19669 27396 19703
rect 27344 19660 27396 19669
rect 27804 19737 27813 19771
rect 27813 19737 27847 19771
rect 27847 19737 27856 19771
rect 27804 19728 27856 19737
rect 29000 19728 29052 19780
rect 31208 19728 31260 19780
rect 31944 19728 31996 19780
rect 34612 19796 34664 19848
rect 38844 20000 38896 20052
rect 40040 20000 40092 20052
rect 40684 20000 40736 20052
rect 42616 20000 42668 20052
rect 41696 19932 41748 19984
rect 43628 20000 43680 20052
rect 50160 20043 50212 20052
rect 35624 19839 35676 19848
rect 35624 19805 35633 19839
rect 35633 19805 35667 19839
rect 35667 19805 35676 19839
rect 35624 19796 35676 19805
rect 38016 19839 38068 19848
rect 38016 19805 38025 19839
rect 38025 19805 38059 19839
rect 38059 19805 38068 19839
rect 38476 19839 38528 19848
rect 38016 19796 38068 19805
rect 38476 19805 38485 19839
rect 38485 19805 38519 19839
rect 38519 19805 38528 19839
rect 38476 19796 38528 19805
rect 27712 19660 27764 19712
rect 31116 19660 31168 19712
rect 32496 19660 32548 19712
rect 36268 19703 36320 19712
rect 36268 19669 36277 19703
rect 36277 19669 36311 19703
rect 36311 19669 36320 19703
rect 36268 19660 36320 19669
rect 38752 19728 38804 19780
rect 39212 19771 39264 19780
rect 39212 19737 39221 19771
rect 39221 19737 39255 19771
rect 39255 19737 39264 19771
rect 39212 19728 39264 19737
rect 38844 19660 38896 19712
rect 40868 19864 40920 19916
rect 41328 19907 41380 19916
rect 41328 19873 41337 19907
rect 41337 19873 41371 19907
rect 41371 19873 41380 19907
rect 41328 19864 41380 19873
rect 41788 19864 41840 19916
rect 43260 19907 43312 19916
rect 43260 19873 43269 19907
rect 43269 19873 43303 19907
rect 43303 19873 43312 19907
rect 43260 19864 43312 19873
rect 50160 20009 50169 20043
rect 50169 20009 50203 20043
rect 50203 20009 50212 20043
rect 50160 20000 50212 20009
rect 50344 20043 50396 20052
rect 50344 20009 50353 20043
rect 50353 20009 50387 20043
rect 50387 20009 50396 20043
rect 50344 20000 50396 20009
rect 50436 20000 50488 20052
rect 53196 20000 53248 20052
rect 52092 19932 52144 19984
rect 52552 19932 52604 19984
rect 53656 19932 53708 19984
rect 42064 19839 42116 19848
rect 42064 19805 42073 19839
rect 42073 19805 42107 19839
rect 42107 19805 42116 19839
rect 42064 19796 42116 19805
rect 43536 19839 43588 19848
rect 43536 19805 43545 19839
rect 43545 19805 43579 19839
rect 43579 19805 43588 19839
rect 43536 19796 43588 19805
rect 44640 19796 44692 19848
rect 39396 19728 39448 19780
rect 45744 19796 45796 19848
rect 50160 19864 50212 19916
rect 52828 19864 52880 19916
rect 53012 19907 53064 19916
rect 53012 19873 53021 19907
rect 53021 19873 53055 19907
rect 53055 19873 53064 19907
rect 53012 19864 53064 19873
rect 50344 19839 50396 19848
rect 42156 19660 42208 19712
rect 44732 19660 44784 19712
rect 46480 19728 46532 19780
rect 48780 19771 48832 19780
rect 48780 19737 48789 19771
rect 48789 19737 48823 19771
rect 48823 19737 48832 19771
rect 48780 19728 48832 19737
rect 49332 19728 49384 19780
rect 50344 19805 50353 19839
rect 50353 19805 50387 19839
rect 50387 19805 50396 19839
rect 50344 19796 50396 19805
rect 50436 19839 50488 19848
rect 50436 19805 50445 19839
rect 50445 19805 50479 19839
rect 50479 19805 50488 19839
rect 51264 19839 51316 19848
rect 50436 19796 50488 19805
rect 51264 19805 51273 19839
rect 51273 19805 51307 19839
rect 51307 19805 51316 19839
rect 51264 19796 51316 19805
rect 52092 19839 52144 19848
rect 50068 19728 50120 19780
rect 50804 19728 50856 19780
rect 46572 19660 46624 19712
rect 48964 19660 49016 19712
rect 51816 19660 51868 19712
rect 52092 19805 52102 19839
rect 52102 19805 52136 19839
rect 52136 19805 52144 19839
rect 52092 19796 52144 19805
rect 53104 19796 53156 19848
rect 53656 19796 53708 19848
rect 53748 19839 53800 19848
rect 53748 19805 53757 19839
rect 53757 19805 53791 19839
rect 53791 19805 53800 19839
rect 53748 19796 53800 19805
rect 54760 19796 54812 19848
rect 55588 19864 55640 19916
rect 56324 19907 56376 19916
rect 56324 19873 56333 19907
rect 56333 19873 56367 19907
rect 56367 19873 56376 19907
rect 56324 19864 56376 19873
rect 53840 19728 53892 19780
rect 52460 19660 52512 19712
rect 53288 19703 53340 19712
rect 53288 19669 53297 19703
rect 53297 19669 53331 19703
rect 53331 19669 53340 19703
rect 53288 19660 53340 19669
rect 57336 19728 57388 19780
rect 15398 19558 15450 19610
rect 15462 19558 15514 19610
rect 15526 19558 15578 19610
rect 15590 19558 15642 19610
rect 15654 19558 15706 19610
rect 29846 19558 29898 19610
rect 29910 19558 29962 19610
rect 29974 19558 30026 19610
rect 30038 19558 30090 19610
rect 30102 19558 30154 19610
rect 44294 19558 44346 19610
rect 44358 19558 44410 19610
rect 44422 19558 44474 19610
rect 44486 19558 44538 19610
rect 44550 19558 44602 19610
rect 6184 19456 6236 19508
rect 4252 19388 4304 19440
rect 5356 19388 5408 19440
rect 7656 19388 7708 19440
rect 9680 19456 9732 19508
rect 11336 19456 11388 19508
rect 12532 19456 12584 19508
rect 14004 19456 14056 19508
rect 14372 19456 14424 19508
rect 17408 19456 17460 19508
rect 18788 19456 18840 19508
rect 19708 19456 19760 19508
rect 2136 19363 2188 19372
rect 2136 19329 2145 19363
rect 2145 19329 2179 19363
rect 2179 19329 2188 19363
rect 2136 19320 2188 19329
rect 6368 19320 6420 19372
rect 7104 19320 7156 19372
rect 10232 19320 10284 19372
rect 10876 19320 10928 19372
rect 11428 19388 11480 19440
rect 12348 19388 12400 19440
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 11888 19320 11940 19372
rect 12992 19363 13044 19372
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 15016 19320 15068 19372
rect 18236 19388 18288 19440
rect 19340 19388 19392 19440
rect 23388 19456 23440 19508
rect 23480 19456 23532 19508
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 3884 19252 3936 19304
rect 4252 19252 4304 19304
rect 6920 19252 6972 19304
rect 5448 19184 5500 19236
rect 9128 19227 9180 19236
rect 9128 19193 9137 19227
rect 9137 19193 9171 19227
rect 9171 19193 9180 19227
rect 9128 19184 9180 19193
rect 12900 19252 12952 19304
rect 13268 19252 13320 19304
rect 17040 19252 17092 19304
rect 17960 19363 18012 19372
rect 17960 19329 17969 19363
rect 17969 19329 18003 19363
rect 18003 19329 18012 19363
rect 17960 19320 18012 19329
rect 18880 19320 18932 19372
rect 19984 19363 20036 19372
rect 19984 19329 19993 19363
rect 19993 19329 20027 19363
rect 20027 19329 20036 19363
rect 19984 19320 20036 19329
rect 22376 19320 22428 19372
rect 25136 19388 25188 19440
rect 24860 19363 24912 19372
rect 24860 19329 24869 19363
rect 24869 19329 24903 19363
rect 24903 19329 24912 19363
rect 24860 19320 24912 19329
rect 27804 19456 27856 19508
rect 31024 19499 31076 19508
rect 31024 19465 31033 19499
rect 31033 19465 31067 19499
rect 31067 19465 31076 19499
rect 31024 19456 31076 19465
rect 27252 19431 27304 19440
rect 27252 19397 27261 19431
rect 27261 19397 27295 19431
rect 27295 19397 27304 19431
rect 27252 19388 27304 19397
rect 30564 19388 30616 19440
rect 19616 19252 19668 19304
rect 16764 19184 16816 19236
rect 19432 19184 19484 19236
rect 25044 19252 25096 19304
rect 23756 19184 23808 19236
rect 31024 19320 31076 19372
rect 36268 19456 36320 19508
rect 40316 19456 40368 19508
rect 42156 19456 42208 19508
rect 43260 19499 43312 19508
rect 43260 19465 43269 19499
rect 43269 19465 43303 19499
rect 43303 19465 43312 19499
rect 43260 19456 43312 19465
rect 48320 19456 48372 19508
rect 51356 19456 51408 19508
rect 53012 19456 53064 19508
rect 53656 19456 53708 19508
rect 35348 19388 35400 19440
rect 41052 19388 41104 19440
rect 29460 19295 29512 19304
rect 29460 19261 29469 19295
rect 29469 19261 29503 19295
rect 29503 19261 29512 19295
rect 29460 19252 29512 19261
rect 30196 19252 30248 19304
rect 34612 19363 34664 19372
rect 34612 19329 34621 19363
rect 34621 19329 34655 19363
rect 34655 19329 34664 19363
rect 34612 19320 34664 19329
rect 35256 19320 35308 19372
rect 37464 19320 37516 19372
rect 39212 19363 39264 19372
rect 39212 19329 39221 19363
rect 39221 19329 39255 19363
rect 39255 19329 39264 19363
rect 39212 19320 39264 19329
rect 41604 19363 41656 19372
rect 41604 19329 41613 19363
rect 41613 19329 41647 19363
rect 41647 19329 41656 19363
rect 41604 19320 41656 19329
rect 42616 19363 42668 19372
rect 42616 19329 42625 19363
rect 42625 19329 42659 19363
rect 42659 19329 42668 19363
rect 42616 19320 42668 19329
rect 43076 19363 43128 19372
rect 43076 19329 43085 19363
rect 43085 19329 43119 19363
rect 43119 19329 43128 19363
rect 43076 19320 43128 19329
rect 46572 19431 46624 19440
rect 43996 19363 44048 19372
rect 43996 19329 44005 19363
rect 44005 19329 44039 19363
rect 44039 19329 44048 19363
rect 44640 19363 44692 19372
rect 43996 19320 44048 19329
rect 44640 19329 44649 19363
rect 44649 19329 44683 19363
rect 44683 19329 44692 19363
rect 44640 19320 44692 19329
rect 45376 19363 45428 19372
rect 45376 19329 45385 19363
rect 45385 19329 45419 19363
rect 45419 19329 45428 19363
rect 45376 19320 45428 19329
rect 46572 19397 46581 19431
rect 46581 19397 46615 19431
rect 46615 19397 46624 19431
rect 46572 19388 46624 19397
rect 45744 19320 45796 19372
rect 46296 19363 46348 19372
rect 26608 19184 26660 19236
rect 32496 19252 32548 19304
rect 35440 19295 35492 19304
rect 35440 19261 35449 19295
rect 35449 19261 35483 19295
rect 35483 19261 35492 19295
rect 35440 19252 35492 19261
rect 36084 19252 36136 19304
rect 38384 19295 38436 19304
rect 35072 19184 35124 19236
rect 38384 19261 38393 19295
rect 38393 19261 38427 19295
rect 38427 19261 38436 19295
rect 38384 19252 38436 19261
rect 46296 19329 46305 19363
rect 46305 19329 46339 19363
rect 46339 19329 46348 19363
rect 46296 19320 46348 19329
rect 47952 19363 48004 19372
rect 47952 19329 47961 19363
rect 47961 19329 47995 19363
rect 47995 19329 48004 19363
rect 47952 19320 48004 19329
rect 48872 19363 48924 19372
rect 48872 19329 48881 19363
rect 48881 19329 48915 19363
rect 48915 19329 48924 19363
rect 48872 19320 48924 19329
rect 50344 19388 50396 19440
rect 50804 19388 50856 19440
rect 51080 19320 51132 19372
rect 51816 19363 51868 19372
rect 51816 19329 51825 19363
rect 51825 19329 51859 19363
rect 51859 19329 51868 19363
rect 51816 19320 51868 19329
rect 52828 19363 52880 19372
rect 52828 19329 52837 19363
rect 52837 19329 52871 19363
rect 52871 19329 52880 19363
rect 52828 19320 52880 19329
rect 53012 19363 53064 19372
rect 53012 19329 53021 19363
rect 53021 19329 53055 19363
rect 53055 19329 53064 19363
rect 53012 19320 53064 19329
rect 46480 19252 46532 19304
rect 47676 19252 47728 19304
rect 48044 19295 48096 19304
rect 48044 19261 48053 19295
rect 48053 19261 48087 19295
rect 48087 19261 48096 19295
rect 48044 19252 48096 19261
rect 48964 19252 49016 19304
rect 49516 19295 49568 19304
rect 49516 19261 49525 19295
rect 49525 19261 49559 19295
rect 49559 19261 49568 19295
rect 49516 19252 49568 19261
rect 51172 19295 51224 19304
rect 51172 19261 51181 19295
rect 51181 19261 51215 19295
rect 51215 19261 51224 19295
rect 51172 19252 51224 19261
rect 57336 19388 57388 19440
rect 53932 19320 53984 19372
rect 54300 19363 54352 19372
rect 54300 19329 54309 19363
rect 54309 19329 54343 19363
rect 54343 19329 54352 19363
rect 54300 19320 54352 19329
rect 52552 19184 52604 19236
rect 53288 19184 53340 19236
rect 3976 19116 4028 19168
rect 9588 19116 9640 19168
rect 11336 19116 11388 19168
rect 13176 19116 13228 19168
rect 17316 19159 17368 19168
rect 17316 19125 17325 19159
rect 17325 19125 17359 19159
rect 17359 19125 17368 19159
rect 17316 19116 17368 19125
rect 21180 19159 21232 19168
rect 21180 19125 21189 19159
rect 21189 19125 21223 19159
rect 21223 19125 21232 19159
rect 21180 19116 21232 19125
rect 24216 19159 24268 19168
rect 24216 19125 24225 19159
rect 24225 19125 24259 19159
rect 24259 19125 24268 19159
rect 24216 19116 24268 19125
rect 26148 19116 26200 19168
rect 30380 19159 30432 19168
rect 30380 19125 30389 19159
rect 30389 19125 30423 19159
rect 30423 19125 30432 19159
rect 30380 19116 30432 19125
rect 33876 19159 33928 19168
rect 33876 19125 33885 19159
rect 33885 19125 33919 19159
rect 33919 19125 33928 19159
rect 33876 19116 33928 19125
rect 44640 19116 44692 19168
rect 46480 19116 46532 19168
rect 51172 19116 51224 19168
rect 53840 19159 53892 19168
rect 53840 19125 53849 19159
rect 53849 19125 53883 19159
rect 53883 19125 53892 19159
rect 53840 19116 53892 19125
rect 8174 19014 8226 19066
rect 8238 19014 8290 19066
rect 8302 19014 8354 19066
rect 8366 19014 8418 19066
rect 8430 19014 8482 19066
rect 22622 19014 22674 19066
rect 22686 19014 22738 19066
rect 22750 19014 22802 19066
rect 22814 19014 22866 19066
rect 22878 19014 22930 19066
rect 37070 19014 37122 19066
rect 37134 19014 37186 19066
rect 37198 19014 37250 19066
rect 37262 19014 37314 19066
rect 37326 19014 37378 19066
rect 51518 19014 51570 19066
rect 51582 19014 51634 19066
rect 51646 19014 51698 19066
rect 51710 19014 51762 19066
rect 51774 19014 51826 19066
rect 11796 18912 11848 18964
rect 2228 18819 2280 18828
rect 2228 18785 2237 18819
rect 2237 18785 2271 18819
rect 2271 18785 2280 18819
rect 2228 18776 2280 18785
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 3056 18708 3108 18760
rect 4252 18751 4304 18760
rect 4252 18717 4261 18751
rect 4261 18717 4295 18751
rect 4295 18717 4304 18751
rect 4252 18708 4304 18717
rect 5908 18751 5960 18760
rect 5908 18717 5917 18751
rect 5917 18717 5951 18751
rect 5951 18717 5960 18751
rect 5908 18708 5960 18717
rect 11336 18844 11388 18896
rect 11520 18844 11572 18896
rect 13360 18776 13412 18828
rect 6644 18683 6696 18692
rect 6644 18649 6653 18683
rect 6653 18649 6687 18683
rect 6687 18649 6696 18683
rect 6644 18640 6696 18649
rect 7104 18640 7156 18692
rect 9864 18640 9916 18692
rect 4896 18615 4948 18624
rect 4896 18581 4905 18615
rect 4905 18581 4939 18615
rect 4939 18581 4948 18615
rect 4896 18572 4948 18581
rect 7288 18572 7340 18624
rect 7472 18572 7524 18624
rect 10232 18615 10284 18624
rect 10232 18581 10241 18615
rect 10241 18581 10275 18615
rect 10275 18581 10284 18615
rect 10232 18572 10284 18581
rect 11336 18572 11388 18624
rect 11520 18615 11572 18624
rect 11520 18581 11529 18615
rect 11529 18581 11563 18615
rect 11563 18581 11572 18615
rect 11520 18572 11572 18581
rect 11888 18708 11940 18760
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 13728 18640 13780 18692
rect 15108 18819 15160 18828
rect 15108 18785 15117 18819
rect 15117 18785 15151 18819
rect 15151 18785 15160 18819
rect 15108 18776 15160 18785
rect 18604 18776 18656 18828
rect 20996 18912 21048 18964
rect 26056 18912 26108 18964
rect 28080 18912 28132 18964
rect 29000 18955 29052 18964
rect 19616 18844 19668 18896
rect 19984 18776 20036 18828
rect 29000 18921 29009 18955
rect 29009 18921 29043 18955
rect 29043 18921 29052 18955
rect 29000 18912 29052 18921
rect 34336 18912 34388 18964
rect 38752 18955 38804 18964
rect 22376 18819 22428 18828
rect 22376 18785 22385 18819
rect 22385 18785 22419 18819
rect 22419 18785 22428 18819
rect 22376 18776 22428 18785
rect 16028 18751 16080 18760
rect 16028 18717 16037 18751
rect 16037 18717 16071 18751
rect 16071 18717 16080 18751
rect 16028 18708 16080 18717
rect 18236 18708 18288 18760
rect 18420 18751 18472 18760
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 17316 18640 17368 18692
rect 13360 18572 13412 18624
rect 14556 18572 14608 18624
rect 17776 18615 17828 18624
rect 17776 18581 17785 18615
rect 17785 18581 17819 18615
rect 17819 18581 17828 18615
rect 17776 18572 17828 18581
rect 18052 18640 18104 18692
rect 20720 18708 20772 18760
rect 21180 18751 21232 18760
rect 21180 18717 21189 18751
rect 21189 18717 21223 18751
rect 21223 18717 21232 18751
rect 22468 18751 22520 18760
rect 21180 18708 21232 18717
rect 22468 18717 22477 18751
rect 22477 18717 22511 18751
rect 22511 18717 22520 18751
rect 22468 18708 22520 18717
rect 23572 18776 23624 18828
rect 29460 18776 29512 18828
rect 23756 18708 23808 18760
rect 24216 18708 24268 18760
rect 25780 18751 25832 18760
rect 25780 18717 25789 18751
rect 25789 18717 25823 18751
rect 25823 18717 25832 18751
rect 25780 18708 25832 18717
rect 25964 18751 26016 18760
rect 25964 18717 25973 18751
rect 25973 18717 26007 18751
rect 26007 18717 26016 18751
rect 25964 18708 26016 18717
rect 30472 18751 30524 18760
rect 30472 18717 30481 18751
rect 30481 18717 30515 18751
rect 30515 18717 30524 18751
rect 30472 18708 30524 18717
rect 31392 18751 31444 18760
rect 31392 18717 31401 18751
rect 31401 18717 31435 18751
rect 31435 18717 31444 18751
rect 38752 18921 38761 18955
rect 38761 18921 38795 18955
rect 38795 18921 38804 18955
rect 38752 18912 38804 18921
rect 36912 18844 36964 18896
rect 45652 18844 45704 18896
rect 40132 18819 40184 18828
rect 31392 18708 31444 18717
rect 21180 18572 21232 18624
rect 21364 18683 21416 18692
rect 21364 18649 21373 18683
rect 21373 18649 21407 18683
rect 21407 18649 21416 18683
rect 21364 18640 21416 18649
rect 26148 18640 26200 18692
rect 27620 18640 27672 18692
rect 27988 18640 28040 18692
rect 32036 18640 32088 18692
rect 33600 18683 33652 18692
rect 33600 18649 33609 18683
rect 33609 18649 33643 18683
rect 33643 18649 33652 18683
rect 33600 18640 33652 18649
rect 33968 18708 34020 18760
rect 36084 18708 36136 18760
rect 40132 18785 40141 18819
rect 40141 18785 40175 18819
rect 40175 18785 40184 18819
rect 40132 18776 40184 18785
rect 43076 18776 43128 18828
rect 49700 18912 49752 18964
rect 49792 18912 49844 18964
rect 50528 18912 50580 18964
rect 52828 18912 52880 18964
rect 53196 18955 53248 18964
rect 53196 18921 53205 18955
rect 53205 18921 53239 18955
rect 53239 18921 53248 18955
rect 53196 18912 53248 18921
rect 52644 18844 52696 18896
rect 48412 18819 48464 18828
rect 48412 18785 48421 18819
rect 48421 18785 48455 18819
rect 48455 18785 48464 18819
rect 48412 18776 48464 18785
rect 34888 18640 34940 18692
rect 24400 18572 24452 18624
rect 26792 18615 26844 18624
rect 26792 18581 26801 18615
rect 26801 18581 26835 18615
rect 26835 18581 26844 18615
rect 26792 18572 26844 18581
rect 29644 18572 29696 18624
rect 36268 18640 36320 18692
rect 39488 18708 39540 18760
rect 41236 18708 41288 18760
rect 42432 18751 42484 18760
rect 42432 18717 42441 18751
rect 42441 18717 42475 18751
rect 42475 18717 42484 18751
rect 42432 18708 42484 18717
rect 43536 18751 43588 18760
rect 43536 18717 43545 18751
rect 43545 18717 43579 18751
rect 43579 18717 43588 18751
rect 43536 18708 43588 18717
rect 43996 18708 44048 18760
rect 44180 18751 44232 18760
rect 44180 18717 44189 18751
rect 44189 18717 44223 18751
rect 44223 18717 44232 18751
rect 44180 18708 44232 18717
rect 46296 18708 46348 18760
rect 47676 18751 47728 18760
rect 47676 18717 47685 18751
rect 47685 18717 47719 18751
rect 47719 18717 47728 18751
rect 47676 18708 47728 18717
rect 48688 18708 48740 18760
rect 50068 18708 50120 18760
rect 52460 18776 52512 18828
rect 52920 18776 52972 18828
rect 53196 18776 53248 18828
rect 54760 18819 54812 18828
rect 54760 18785 54769 18819
rect 54769 18785 54803 18819
rect 54803 18785 54812 18819
rect 54760 18776 54812 18785
rect 41420 18572 41472 18624
rect 41604 18615 41656 18624
rect 41604 18581 41613 18615
rect 41613 18581 41647 18615
rect 41647 18581 41656 18615
rect 41604 18572 41656 18581
rect 42800 18572 42852 18624
rect 44640 18640 44692 18692
rect 45928 18640 45980 18692
rect 47400 18640 47452 18692
rect 52184 18708 52236 18760
rect 57336 18708 57388 18760
rect 50804 18640 50856 18692
rect 52368 18640 52420 18692
rect 57428 18640 57480 18692
rect 51172 18572 51224 18624
rect 54208 18572 54260 18624
rect 15398 18470 15450 18522
rect 15462 18470 15514 18522
rect 15526 18470 15578 18522
rect 15590 18470 15642 18522
rect 15654 18470 15706 18522
rect 29846 18470 29898 18522
rect 29910 18470 29962 18522
rect 29974 18470 30026 18522
rect 30038 18470 30090 18522
rect 30102 18470 30154 18522
rect 44294 18470 44346 18522
rect 44358 18470 44410 18522
rect 44422 18470 44474 18522
rect 44486 18470 44538 18522
rect 44550 18470 44602 18522
rect 4344 18368 4396 18420
rect 5080 18411 5132 18420
rect 5080 18377 5089 18411
rect 5089 18377 5123 18411
rect 5123 18377 5132 18411
rect 5080 18368 5132 18377
rect 6276 18368 6328 18420
rect 7012 18368 7064 18420
rect 10232 18368 10284 18420
rect 11244 18368 11296 18420
rect 14648 18411 14700 18420
rect 14648 18377 14657 18411
rect 14657 18377 14691 18411
rect 14691 18377 14700 18411
rect 14648 18368 14700 18377
rect 16488 18368 16540 18420
rect 19524 18368 19576 18420
rect 21180 18411 21232 18420
rect 21180 18377 21189 18411
rect 21189 18377 21223 18411
rect 21223 18377 21232 18411
rect 21180 18368 21232 18377
rect 22100 18368 22152 18420
rect 4712 18300 4764 18352
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 4068 18232 4120 18284
rect 5632 18275 5684 18284
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 3792 18164 3844 18216
rect 3976 18207 4028 18216
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 5632 18241 5641 18275
rect 5641 18241 5675 18275
rect 5675 18241 5684 18275
rect 5632 18232 5684 18241
rect 5908 18232 5960 18284
rect 6276 18164 6328 18216
rect 6460 18071 6512 18080
rect 6460 18037 6469 18071
rect 6469 18037 6503 18071
rect 6503 18037 6512 18071
rect 6460 18028 6512 18037
rect 7288 18300 7340 18352
rect 13084 18300 13136 18352
rect 13268 18300 13320 18352
rect 11704 18232 11756 18284
rect 13176 18275 13228 18284
rect 11336 18164 11388 18216
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 18420 18300 18472 18352
rect 18696 18300 18748 18352
rect 24860 18368 24912 18420
rect 25044 18368 25096 18420
rect 29644 18368 29696 18420
rect 30196 18368 30248 18420
rect 33968 18368 34020 18420
rect 34888 18368 34940 18420
rect 18972 18275 19024 18284
rect 18972 18241 18981 18275
rect 18981 18241 19015 18275
rect 19015 18241 19024 18275
rect 18972 18232 19024 18241
rect 19064 18232 19116 18284
rect 18696 18164 18748 18216
rect 22100 18232 22152 18284
rect 24952 18300 25004 18352
rect 25688 18300 25740 18352
rect 26056 18300 26108 18352
rect 30656 18300 30708 18352
rect 31944 18300 31996 18352
rect 24676 18207 24728 18216
rect 24676 18173 24685 18207
rect 24685 18173 24719 18207
rect 24719 18173 24728 18207
rect 24676 18164 24728 18173
rect 25228 18164 25280 18216
rect 26148 18207 26200 18216
rect 26148 18173 26157 18207
rect 26157 18173 26191 18207
rect 26191 18173 26200 18207
rect 26148 18164 26200 18173
rect 27436 18232 27488 18284
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 27712 18164 27764 18216
rect 28080 18164 28132 18216
rect 11980 18096 12032 18148
rect 16028 18139 16080 18148
rect 16028 18105 16037 18139
rect 16037 18105 16071 18139
rect 16071 18105 16080 18139
rect 16028 18096 16080 18105
rect 21824 18096 21876 18148
rect 26240 18096 26292 18148
rect 30472 18232 30524 18284
rect 30932 18275 30984 18284
rect 30932 18241 30941 18275
rect 30941 18241 30975 18275
rect 30975 18241 30984 18275
rect 30932 18232 30984 18241
rect 31116 18232 31168 18284
rect 31208 18232 31260 18284
rect 33876 18300 33928 18352
rect 32588 18275 32640 18284
rect 32588 18241 32597 18275
rect 32597 18241 32631 18275
rect 32631 18241 32640 18275
rect 32588 18232 32640 18241
rect 33140 18232 33192 18284
rect 35164 18300 35216 18352
rect 35440 18368 35492 18420
rect 41052 18411 41104 18420
rect 36544 18300 36596 18352
rect 38384 18300 38436 18352
rect 41052 18377 41061 18411
rect 41061 18377 41095 18411
rect 41095 18377 41104 18411
rect 41052 18368 41104 18377
rect 48780 18368 48832 18420
rect 42064 18300 42116 18352
rect 29276 18207 29328 18216
rect 29276 18173 29285 18207
rect 29285 18173 29319 18207
rect 29319 18173 29328 18207
rect 29276 18164 29328 18173
rect 34244 18164 34296 18216
rect 34612 18207 34664 18216
rect 34612 18173 34621 18207
rect 34621 18173 34655 18207
rect 34655 18173 34664 18207
rect 34612 18164 34664 18173
rect 34796 18164 34848 18216
rect 36452 18164 36504 18216
rect 38476 18232 38528 18284
rect 40868 18232 40920 18284
rect 41696 18232 41748 18284
rect 42524 18300 42576 18352
rect 42616 18232 42668 18284
rect 43352 18275 43404 18284
rect 43352 18241 43361 18275
rect 43361 18241 43395 18275
rect 43395 18241 43404 18275
rect 43352 18232 43404 18241
rect 44640 18300 44692 18352
rect 45560 18300 45612 18352
rect 45836 18300 45888 18352
rect 49608 18368 49660 18420
rect 50252 18300 50304 18352
rect 52736 18300 52788 18352
rect 50804 18275 50856 18284
rect 50804 18241 50813 18275
rect 50813 18241 50847 18275
rect 50847 18241 50856 18275
rect 50804 18232 50856 18241
rect 51080 18232 51132 18284
rect 52000 18275 52052 18284
rect 38108 18207 38160 18216
rect 38108 18173 38117 18207
rect 38117 18173 38151 18207
rect 38151 18173 38160 18207
rect 38108 18164 38160 18173
rect 34704 18096 34756 18148
rect 8576 18028 8628 18080
rect 9220 18028 9272 18080
rect 11612 18071 11664 18080
rect 11612 18037 11621 18071
rect 11621 18037 11655 18071
rect 11655 18037 11664 18071
rect 11612 18028 11664 18037
rect 14096 18071 14148 18080
rect 14096 18037 14105 18071
rect 14105 18037 14139 18071
rect 14139 18037 14148 18071
rect 14096 18028 14148 18037
rect 20260 18071 20312 18080
rect 20260 18037 20269 18071
rect 20269 18037 20303 18071
rect 20303 18037 20312 18071
rect 20260 18028 20312 18037
rect 21180 18028 21232 18080
rect 22468 18028 22520 18080
rect 33232 18071 33284 18080
rect 33232 18037 33241 18071
rect 33241 18037 33275 18071
rect 33275 18037 33284 18071
rect 33232 18028 33284 18037
rect 33968 18071 34020 18080
rect 33968 18037 33977 18071
rect 33977 18037 34011 18071
rect 34011 18037 34020 18071
rect 33968 18028 34020 18037
rect 34244 18028 34296 18080
rect 39488 18028 39540 18080
rect 41420 18164 41472 18216
rect 42340 18164 42392 18216
rect 45928 18207 45980 18216
rect 42432 18096 42484 18148
rect 43812 18096 43864 18148
rect 45928 18173 45937 18207
rect 45937 18173 45971 18207
rect 45971 18173 45980 18207
rect 45928 18164 45980 18173
rect 46848 18207 46900 18216
rect 46848 18173 46857 18207
rect 46857 18173 46891 18207
rect 46891 18173 46900 18207
rect 46848 18164 46900 18173
rect 47032 18207 47084 18216
rect 47032 18173 47041 18207
rect 47041 18173 47075 18207
rect 47075 18173 47084 18207
rect 47032 18164 47084 18173
rect 46756 18096 46808 18148
rect 48596 18096 48648 18148
rect 41420 18028 41472 18080
rect 42984 18028 43036 18080
rect 43996 18028 44048 18080
rect 50068 18164 50120 18216
rect 50528 18207 50580 18216
rect 50528 18173 50537 18207
rect 50537 18173 50571 18207
rect 50571 18173 50580 18207
rect 50528 18164 50580 18173
rect 52000 18241 52009 18275
rect 52009 18241 52043 18275
rect 52043 18241 52052 18275
rect 52000 18232 52052 18241
rect 52184 18275 52236 18284
rect 52184 18241 52193 18275
rect 52193 18241 52227 18275
rect 52227 18241 52236 18275
rect 52184 18232 52236 18241
rect 52828 18232 52880 18284
rect 53288 18232 53340 18284
rect 56416 18232 56468 18284
rect 57888 18275 57940 18284
rect 57888 18241 57897 18275
rect 57897 18241 57931 18275
rect 57931 18241 57940 18275
rect 57888 18232 57940 18241
rect 53012 18096 53064 18148
rect 53196 18207 53248 18216
rect 53196 18173 53205 18207
rect 53205 18173 53239 18207
rect 53239 18173 53248 18207
rect 53196 18164 53248 18173
rect 54116 18164 54168 18216
rect 56232 18207 56284 18216
rect 56232 18173 56241 18207
rect 56241 18173 56275 18207
rect 56275 18173 56284 18207
rect 56232 18164 56284 18173
rect 53472 18096 53524 18148
rect 56692 18139 56744 18148
rect 56692 18105 56701 18139
rect 56701 18105 56735 18139
rect 56735 18105 56744 18139
rect 56692 18096 56744 18105
rect 49056 18071 49108 18080
rect 49056 18037 49065 18071
rect 49065 18037 49099 18071
rect 49099 18037 49108 18071
rect 49056 18028 49108 18037
rect 50436 18028 50488 18080
rect 53564 18028 53616 18080
rect 53840 18071 53892 18080
rect 53840 18037 53849 18071
rect 53849 18037 53883 18071
rect 53883 18037 53892 18071
rect 53840 18028 53892 18037
rect 55956 18028 56008 18080
rect 57796 18028 57848 18080
rect 8174 17926 8226 17978
rect 8238 17926 8290 17978
rect 8302 17926 8354 17978
rect 8366 17926 8418 17978
rect 8430 17926 8482 17978
rect 22622 17926 22674 17978
rect 22686 17926 22738 17978
rect 22750 17926 22802 17978
rect 22814 17926 22866 17978
rect 22878 17926 22930 17978
rect 37070 17926 37122 17978
rect 37134 17926 37186 17978
rect 37198 17926 37250 17978
rect 37262 17926 37314 17978
rect 37326 17926 37378 17978
rect 51518 17926 51570 17978
rect 51582 17926 51634 17978
rect 51646 17926 51698 17978
rect 51710 17926 51762 17978
rect 51774 17926 51826 17978
rect 2136 17824 2188 17876
rect 11060 17824 11112 17876
rect 11428 17824 11480 17876
rect 15292 17824 15344 17876
rect 16212 17824 16264 17876
rect 20260 17824 20312 17876
rect 22928 17824 22980 17876
rect 23020 17824 23072 17876
rect 23572 17824 23624 17876
rect 24952 17824 25004 17876
rect 36820 17824 36872 17876
rect 38292 17867 38344 17876
rect 38292 17833 38301 17867
rect 38301 17833 38335 17867
rect 38335 17833 38344 17867
rect 38292 17824 38344 17833
rect 41420 17824 41472 17876
rect 41880 17824 41932 17876
rect 42524 17824 42576 17876
rect 50528 17824 50580 17876
rect 2872 17688 2924 17740
rect 3056 17620 3108 17672
rect 4252 17756 4304 17808
rect 5172 17688 5224 17740
rect 11520 17756 11572 17808
rect 11888 17756 11940 17808
rect 18604 17799 18656 17808
rect 18604 17765 18613 17799
rect 18613 17765 18647 17799
rect 18647 17765 18656 17799
rect 18604 17756 18656 17765
rect 18696 17756 18748 17808
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 5632 17620 5684 17672
rect 9588 17663 9640 17672
rect 5724 17595 5776 17604
rect 5724 17561 5733 17595
rect 5733 17561 5767 17595
rect 5767 17561 5776 17595
rect 5724 17552 5776 17561
rect 9588 17629 9597 17663
rect 9597 17629 9631 17663
rect 9631 17629 9640 17663
rect 9588 17620 9640 17629
rect 15936 17731 15988 17740
rect 15936 17697 15945 17731
rect 15945 17697 15979 17731
rect 15979 17697 15988 17731
rect 15936 17688 15988 17697
rect 11704 17620 11756 17672
rect 15200 17620 15252 17672
rect 6828 17552 6880 17604
rect 1952 17484 2004 17536
rect 6460 17484 6512 17536
rect 8668 17484 8720 17536
rect 9772 17552 9824 17604
rect 11796 17595 11848 17604
rect 11796 17561 11805 17595
rect 11805 17561 11839 17595
rect 11839 17561 11848 17595
rect 11796 17552 11848 17561
rect 18420 17552 18472 17604
rect 19800 17620 19852 17672
rect 20444 17663 20496 17672
rect 19340 17552 19392 17604
rect 20444 17629 20453 17663
rect 20453 17629 20487 17663
rect 20487 17629 20496 17663
rect 20444 17620 20496 17629
rect 20628 17620 20680 17672
rect 20996 17552 21048 17604
rect 11888 17484 11940 17536
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 17592 17484 17644 17536
rect 20444 17484 20496 17536
rect 22376 17620 22428 17672
rect 24676 17756 24728 17808
rect 30564 17756 30616 17808
rect 31576 17756 31628 17808
rect 25964 17620 26016 17672
rect 26148 17620 26200 17672
rect 28724 17688 28776 17740
rect 37188 17756 37240 17808
rect 42892 17756 42944 17808
rect 52184 17824 52236 17876
rect 53196 17824 53248 17876
rect 53932 17867 53984 17876
rect 53932 17833 53941 17867
rect 53941 17833 53975 17867
rect 53975 17833 53984 17867
rect 53932 17824 53984 17833
rect 56416 17824 56468 17876
rect 32036 17688 32088 17740
rect 34796 17688 34848 17740
rect 36268 17688 36320 17740
rect 38936 17688 38988 17740
rect 41604 17688 41656 17740
rect 43812 17731 43864 17740
rect 43812 17697 43821 17731
rect 43821 17697 43855 17731
rect 43855 17697 43864 17731
rect 43812 17688 43864 17697
rect 47400 17688 47452 17740
rect 47676 17688 47728 17740
rect 48044 17688 48096 17740
rect 31668 17620 31720 17672
rect 35256 17663 35308 17672
rect 35256 17629 35265 17663
rect 35265 17629 35299 17663
rect 35299 17629 35308 17663
rect 35256 17620 35308 17629
rect 35900 17663 35952 17672
rect 35900 17629 35909 17663
rect 35909 17629 35943 17663
rect 35943 17629 35952 17663
rect 35900 17620 35952 17629
rect 38108 17663 38160 17672
rect 38108 17629 38117 17663
rect 38117 17629 38151 17663
rect 38151 17629 38160 17663
rect 38108 17620 38160 17629
rect 40316 17663 40368 17672
rect 40316 17629 40325 17663
rect 40325 17629 40359 17663
rect 40359 17629 40368 17663
rect 40316 17620 40368 17629
rect 23848 17552 23900 17604
rect 27344 17552 27396 17604
rect 31208 17595 31260 17604
rect 29736 17484 29788 17536
rect 31208 17561 31217 17595
rect 31217 17561 31251 17595
rect 31251 17561 31260 17595
rect 31208 17552 31260 17561
rect 32312 17552 32364 17604
rect 35808 17552 35860 17604
rect 36176 17595 36228 17604
rect 36176 17561 36185 17595
rect 36185 17561 36219 17595
rect 36219 17561 36228 17595
rect 36176 17552 36228 17561
rect 33324 17484 33376 17536
rect 34060 17527 34112 17536
rect 34060 17493 34069 17527
rect 34069 17493 34103 17527
rect 34103 17493 34112 17527
rect 34060 17484 34112 17493
rect 34612 17484 34664 17536
rect 38844 17552 38896 17604
rect 39120 17595 39172 17604
rect 39120 17561 39129 17595
rect 39129 17561 39163 17595
rect 39163 17561 39172 17595
rect 39120 17552 39172 17561
rect 41236 17620 41288 17672
rect 42064 17620 42116 17672
rect 44180 17663 44232 17672
rect 44180 17629 44189 17663
rect 44189 17629 44223 17663
rect 44223 17629 44232 17663
rect 44180 17620 44232 17629
rect 45008 17663 45060 17672
rect 45008 17629 45017 17663
rect 45017 17629 45051 17663
rect 45051 17629 45060 17663
rect 45008 17620 45060 17629
rect 50436 17731 50488 17740
rect 50436 17697 50445 17731
rect 50445 17697 50479 17731
rect 50479 17697 50488 17731
rect 50436 17688 50488 17697
rect 48320 17663 48372 17672
rect 48320 17629 48329 17663
rect 48329 17629 48363 17663
rect 48363 17629 48372 17663
rect 48320 17620 48372 17629
rect 49056 17620 49108 17672
rect 52368 17688 52420 17740
rect 51816 17663 51868 17672
rect 38292 17484 38344 17536
rect 40960 17484 41012 17536
rect 41788 17484 41840 17536
rect 42800 17552 42852 17604
rect 45192 17595 45244 17604
rect 45192 17561 45201 17595
rect 45201 17561 45235 17595
rect 45235 17561 45244 17595
rect 45192 17552 45244 17561
rect 45928 17552 45980 17604
rect 49516 17484 49568 17536
rect 51816 17629 51825 17663
rect 51825 17629 51859 17663
rect 51859 17629 51868 17663
rect 51816 17620 51868 17629
rect 52460 17663 52512 17672
rect 52184 17552 52236 17604
rect 52460 17629 52469 17663
rect 52469 17629 52503 17663
rect 52503 17629 52512 17663
rect 52460 17620 52512 17629
rect 52920 17663 52972 17672
rect 52920 17629 52929 17663
rect 52929 17629 52963 17663
rect 52963 17629 52972 17663
rect 52920 17620 52972 17629
rect 54300 17688 54352 17740
rect 56324 17688 56376 17740
rect 56692 17731 56744 17740
rect 56692 17697 56701 17731
rect 56701 17697 56735 17731
rect 56735 17697 56744 17731
rect 56692 17688 56744 17697
rect 54116 17663 54168 17672
rect 52736 17552 52788 17604
rect 53012 17484 53064 17536
rect 54116 17629 54125 17663
rect 54125 17629 54159 17663
rect 54159 17629 54168 17663
rect 54116 17620 54168 17629
rect 54760 17620 54812 17672
rect 53472 17595 53524 17604
rect 53472 17561 53481 17595
rect 53481 17561 53515 17595
rect 53515 17561 53524 17595
rect 53472 17552 53524 17561
rect 53288 17527 53340 17536
rect 53288 17493 53297 17527
rect 53297 17493 53331 17527
rect 53331 17493 53340 17527
rect 54392 17595 54444 17604
rect 54392 17561 54401 17595
rect 54401 17561 54435 17595
rect 54435 17561 54444 17595
rect 54392 17552 54444 17561
rect 56784 17552 56836 17604
rect 57336 17552 57388 17604
rect 53288 17484 53340 17493
rect 56692 17484 56744 17536
rect 15398 17382 15450 17434
rect 15462 17382 15514 17434
rect 15526 17382 15578 17434
rect 15590 17382 15642 17434
rect 15654 17382 15706 17434
rect 29846 17382 29898 17434
rect 29910 17382 29962 17434
rect 29974 17382 30026 17434
rect 30038 17382 30090 17434
rect 30102 17382 30154 17434
rect 44294 17382 44346 17434
rect 44358 17382 44410 17434
rect 44422 17382 44474 17434
rect 44486 17382 44538 17434
rect 44550 17382 44602 17434
rect 5356 17280 5408 17332
rect 7012 17280 7064 17332
rect 8576 17280 8628 17332
rect 17592 17280 17644 17332
rect 1952 17255 2004 17264
rect 1952 17221 1961 17255
rect 1961 17221 1995 17255
rect 1995 17221 2004 17255
rect 1952 17212 2004 17221
rect 3516 17212 3568 17264
rect 4804 17212 4856 17264
rect 11612 17212 11664 17264
rect 15292 17212 15344 17264
rect 17960 17212 18012 17264
rect 19800 17280 19852 17332
rect 25044 17323 25096 17332
rect 25044 17289 25053 17323
rect 25053 17289 25087 17323
rect 25087 17289 25096 17323
rect 25044 17280 25096 17289
rect 25688 17323 25740 17332
rect 25688 17289 25697 17323
rect 25697 17289 25731 17323
rect 25731 17289 25740 17323
rect 25688 17280 25740 17289
rect 22928 17212 22980 17264
rect 3056 17008 3108 17060
rect 5908 17144 5960 17196
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 9128 17144 9180 17196
rect 10324 17187 10376 17196
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 10784 17187 10836 17196
rect 10784 17153 10793 17187
rect 10793 17153 10827 17187
rect 10827 17153 10836 17187
rect 10784 17144 10836 17153
rect 16488 17144 16540 17196
rect 5448 17076 5500 17128
rect 6736 17076 6788 17128
rect 5264 17008 5316 17060
rect 8760 17076 8812 17128
rect 11060 17076 11112 17128
rect 16580 17076 16632 17128
rect 17960 17076 18012 17128
rect 20720 17119 20772 17128
rect 20720 17085 20729 17119
rect 20729 17085 20763 17119
rect 20763 17085 20772 17119
rect 20720 17076 20772 17085
rect 7380 17008 7432 17060
rect 12256 17008 12308 17060
rect 21180 17051 21232 17060
rect 21180 17017 21189 17051
rect 21189 17017 21223 17051
rect 21223 17017 21232 17051
rect 21180 17008 21232 17017
rect 21824 17185 21876 17196
rect 21824 17151 21833 17185
rect 21833 17151 21867 17185
rect 21867 17151 21876 17185
rect 21824 17144 21876 17151
rect 23296 17187 23348 17196
rect 23296 17153 23305 17187
rect 23305 17153 23339 17187
rect 23339 17153 23348 17187
rect 23296 17144 23348 17153
rect 24860 17144 24912 17196
rect 28080 17144 28132 17196
rect 28356 17187 28408 17196
rect 28356 17153 28365 17187
rect 28365 17153 28399 17187
rect 28399 17153 28408 17187
rect 28356 17144 28408 17153
rect 31392 17144 31444 17196
rect 24952 17076 25004 17128
rect 29184 17119 29236 17128
rect 29184 17085 29193 17119
rect 29193 17085 29227 17119
rect 29227 17085 29236 17119
rect 29184 17076 29236 17085
rect 29276 17076 29328 17128
rect 30104 17076 30156 17128
rect 32588 17212 32640 17264
rect 34796 17212 34848 17264
rect 34704 17187 34756 17196
rect 34704 17153 34713 17187
rect 34713 17153 34747 17187
rect 34747 17153 34756 17187
rect 34704 17144 34756 17153
rect 37188 17280 37240 17332
rect 35808 17212 35860 17264
rect 38568 17280 38620 17332
rect 44180 17280 44232 17332
rect 44824 17280 44876 17332
rect 38844 17212 38896 17264
rect 40776 17212 40828 17264
rect 46756 17280 46808 17332
rect 48596 17323 48648 17332
rect 48596 17289 48605 17323
rect 48605 17289 48639 17323
rect 48639 17289 48648 17323
rect 48596 17280 48648 17289
rect 51816 17280 51868 17332
rect 53472 17280 53524 17332
rect 53564 17280 53616 17332
rect 56232 17280 56284 17332
rect 57888 17323 57940 17332
rect 57888 17289 57897 17323
rect 57897 17289 57931 17323
rect 57931 17289 57940 17323
rect 57888 17280 57940 17289
rect 36452 17144 36504 17196
rect 39488 17187 39540 17196
rect 39488 17153 39497 17187
rect 39497 17153 39531 17187
rect 39531 17153 39540 17187
rect 39488 17144 39540 17153
rect 41788 17144 41840 17196
rect 32220 17119 32272 17128
rect 32220 17085 32229 17119
rect 32229 17085 32263 17119
rect 32263 17085 32272 17119
rect 32220 17076 32272 17085
rect 33232 17076 33284 17128
rect 35992 17076 36044 17128
rect 38568 17076 38620 17128
rect 39764 17119 39816 17128
rect 39764 17085 39773 17119
rect 39773 17085 39807 17119
rect 39807 17085 39816 17119
rect 39764 17076 39816 17085
rect 28816 17008 28868 17060
rect 29644 17051 29696 17060
rect 29644 17017 29653 17051
rect 29653 17017 29687 17051
rect 29687 17017 29696 17051
rect 29644 17008 29696 17017
rect 3148 16940 3200 16992
rect 3424 16940 3476 16992
rect 12716 16940 12768 16992
rect 18236 16940 18288 16992
rect 22284 16940 22336 16992
rect 23204 16940 23256 16992
rect 25044 16940 25096 16992
rect 26424 16940 26476 16992
rect 26976 16983 27028 16992
rect 26976 16949 26985 16983
rect 26985 16949 27019 16983
rect 27019 16949 27028 16983
rect 26976 16940 27028 16949
rect 31024 16940 31076 16992
rect 31300 16983 31352 16992
rect 31300 16949 31309 16983
rect 31309 16949 31343 16983
rect 31343 16949 31352 16983
rect 31300 16940 31352 16949
rect 32588 16940 32640 16992
rect 36360 17008 36412 17060
rect 42892 17076 42944 17128
rect 43536 17008 43588 17060
rect 45652 17076 45704 17128
rect 45928 17119 45980 17128
rect 45928 17085 45937 17119
rect 45937 17085 45971 17119
rect 45971 17085 45980 17119
rect 45928 17076 45980 17085
rect 49056 17212 49108 17264
rect 47768 17187 47820 17196
rect 47768 17153 47777 17187
rect 47777 17153 47811 17187
rect 47811 17153 47820 17187
rect 47768 17144 47820 17153
rect 48044 17187 48096 17196
rect 48044 17153 48053 17187
rect 48053 17153 48087 17187
rect 48087 17153 48096 17187
rect 48044 17144 48096 17153
rect 49792 17212 49844 17264
rect 50252 17212 50304 17264
rect 52920 17255 52972 17264
rect 52920 17221 52929 17255
rect 52929 17221 52963 17255
rect 52963 17221 52972 17255
rect 55956 17255 56008 17264
rect 52920 17212 52972 17221
rect 55956 17221 55965 17255
rect 55965 17221 55999 17255
rect 55999 17221 56008 17255
rect 55956 17212 56008 17221
rect 48136 17008 48188 17060
rect 36084 16983 36136 16992
rect 36084 16949 36093 16983
rect 36093 16949 36127 16983
rect 36127 16949 36136 16983
rect 36084 16940 36136 16949
rect 38292 16940 38344 16992
rect 39028 16983 39080 16992
rect 39028 16949 39037 16983
rect 39037 16949 39071 16983
rect 39071 16949 39080 16983
rect 39028 16940 39080 16949
rect 41236 16983 41288 16992
rect 41236 16949 41245 16983
rect 41245 16949 41279 16983
rect 41279 16949 41288 16983
rect 41236 16940 41288 16949
rect 47676 16940 47728 16992
rect 51908 17187 51960 17196
rect 51908 17153 51917 17187
rect 51917 17153 51951 17187
rect 51951 17153 51960 17187
rect 51908 17144 51960 17153
rect 52552 17144 52604 17196
rect 52736 17187 52788 17196
rect 52736 17153 52745 17187
rect 52745 17153 52779 17187
rect 52779 17153 52788 17187
rect 52736 17144 52788 17153
rect 55036 17187 55088 17196
rect 55036 17153 55045 17187
rect 55045 17153 55079 17187
rect 55079 17153 55088 17187
rect 55036 17144 55088 17153
rect 55220 17144 55272 17196
rect 50160 17076 50212 17128
rect 52368 17076 52420 17128
rect 54208 17119 54260 17128
rect 54208 17085 54217 17119
rect 54217 17085 54251 17119
rect 54251 17085 54260 17119
rect 54208 17076 54260 17085
rect 51448 17008 51500 17060
rect 51356 16940 51408 16992
rect 52184 17008 52236 17060
rect 53932 17008 53984 17060
rect 57244 17051 57296 17060
rect 57244 17017 57253 17051
rect 57253 17017 57287 17051
rect 57287 17017 57296 17051
rect 57244 17008 57296 17017
rect 52552 16940 52604 16992
rect 52736 16940 52788 16992
rect 53196 16940 53248 16992
rect 8174 16838 8226 16890
rect 8238 16838 8290 16890
rect 8302 16838 8354 16890
rect 8366 16838 8418 16890
rect 8430 16838 8482 16890
rect 22622 16838 22674 16890
rect 22686 16838 22738 16890
rect 22750 16838 22802 16890
rect 22814 16838 22866 16890
rect 22878 16838 22930 16890
rect 37070 16838 37122 16890
rect 37134 16838 37186 16890
rect 37198 16838 37250 16890
rect 37262 16838 37314 16890
rect 37326 16838 37378 16890
rect 51518 16838 51570 16890
rect 51582 16838 51634 16890
rect 51646 16838 51698 16890
rect 51710 16838 51762 16890
rect 51774 16838 51826 16890
rect 3884 16575 3936 16584
rect 3884 16541 3893 16575
rect 3893 16541 3927 16575
rect 3927 16541 3936 16575
rect 3884 16532 3936 16541
rect 6092 16736 6144 16788
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 6552 16600 6604 16652
rect 9036 16668 9088 16720
rect 16580 16736 16632 16788
rect 17776 16736 17828 16788
rect 17868 16736 17920 16788
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 5172 16532 5224 16541
rect 5448 16532 5500 16584
rect 7196 16532 7248 16584
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 10784 16600 10836 16652
rect 5356 16464 5408 16516
rect 5540 16464 5592 16516
rect 6368 16464 6420 16516
rect 8760 16532 8812 16584
rect 9220 16575 9272 16584
rect 9220 16541 9229 16575
rect 9229 16541 9263 16575
rect 9263 16541 9272 16575
rect 9220 16532 9272 16541
rect 11244 16600 11296 16652
rect 13268 16668 13320 16720
rect 16488 16668 16540 16720
rect 14832 16600 14884 16652
rect 15016 16600 15068 16652
rect 16580 16600 16632 16652
rect 19340 16668 19392 16720
rect 23020 16736 23072 16788
rect 24676 16736 24728 16788
rect 25780 16736 25832 16788
rect 18236 16600 18288 16652
rect 20812 16643 20864 16652
rect 4712 16396 4764 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 11336 16396 11388 16448
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 17868 16575 17920 16584
rect 17868 16541 17877 16575
rect 17877 16541 17911 16575
rect 17911 16541 17920 16575
rect 20812 16609 20821 16643
rect 20821 16609 20855 16643
rect 20855 16609 20864 16643
rect 20812 16600 20864 16609
rect 21088 16643 21140 16652
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 21180 16600 21232 16652
rect 17868 16532 17920 16541
rect 18420 16575 18472 16584
rect 18420 16541 18429 16575
rect 18429 16541 18463 16575
rect 18463 16541 18472 16575
rect 25412 16600 25464 16652
rect 25964 16668 26016 16720
rect 30104 16736 30156 16788
rect 29552 16643 29604 16652
rect 18420 16532 18472 16541
rect 23480 16532 23532 16584
rect 29552 16609 29561 16643
rect 29561 16609 29595 16643
rect 29595 16609 29604 16643
rect 29552 16600 29604 16609
rect 33140 16736 33192 16788
rect 33324 16779 33376 16788
rect 33324 16745 33333 16779
rect 33333 16745 33367 16779
rect 33367 16745 33376 16779
rect 33324 16736 33376 16745
rect 35900 16736 35952 16788
rect 39764 16736 39816 16788
rect 40776 16736 40828 16788
rect 42800 16736 42852 16788
rect 44088 16736 44140 16788
rect 44272 16736 44324 16788
rect 47032 16736 47084 16788
rect 35808 16668 35860 16720
rect 31300 16643 31352 16652
rect 31300 16609 31309 16643
rect 31309 16609 31343 16643
rect 31343 16609 31352 16643
rect 31300 16600 31352 16609
rect 33968 16600 34020 16652
rect 41788 16668 41840 16720
rect 43168 16668 43220 16720
rect 36360 16643 36412 16652
rect 27712 16532 27764 16584
rect 28172 16532 28224 16584
rect 29736 16532 29788 16584
rect 31024 16575 31076 16584
rect 18604 16464 18656 16516
rect 22284 16464 22336 16516
rect 15200 16396 15252 16448
rect 15752 16396 15804 16448
rect 16120 16439 16172 16448
rect 16120 16405 16129 16439
rect 16129 16405 16163 16439
rect 16163 16405 16172 16439
rect 16120 16396 16172 16405
rect 16304 16396 16356 16448
rect 20996 16396 21048 16448
rect 24676 16396 24728 16448
rect 27620 16396 27672 16448
rect 28632 16439 28684 16448
rect 28632 16405 28641 16439
rect 28641 16405 28675 16439
rect 28675 16405 28684 16439
rect 28632 16396 28684 16405
rect 28816 16439 28868 16448
rect 28816 16405 28825 16439
rect 28825 16405 28859 16439
rect 28859 16405 28868 16439
rect 28816 16396 28868 16405
rect 31024 16541 31033 16575
rect 31033 16541 31067 16575
rect 31067 16541 31076 16575
rect 31024 16532 31076 16541
rect 36360 16609 36369 16643
rect 36369 16609 36403 16643
rect 36403 16609 36412 16643
rect 36360 16600 36412 16609
rect 37648 16600 37700 16652
rect 38292 16600 38344 16652
rect 34796 16575 34848 16584
rect 34796 16541 34805 16575
rect 34805 16541 34839 16575
rect 34839 16541 34848 16575
rect 34796 16532 34848 16541
rect 31760 16464 31812 16516
rect 34244 16464 34296 16516
rect 35348 16532 35400 16584
rect 35532 16575 35584 16584
rect 35532 16541 35541 16575
rect 35541 16541 35575 16575
rect 35575 16541 35584 16575
rect 40684 16600 40736 16652
rect 42616 16643 42668 16652
rect 42616 16609 42625 16643
rect 42625 16609 42659 16643
rect 42659 16609 42668 16643
rect 42616 16600 42668 16609
rect 44916 16668 44968 16720
rect 44180 16600 44232 16652
rect 35532 16532 35584 16541
rect 44640 16600 44692 16652
rect 33876 16396 33928 16448
rect 34060 16439 34112 16448
rect 34060 16405 34069 16439
rect 34069 16405 34103 16439
rect 34103 16405 34112 16439
rect 34060 16396 34112 16405
rect 41512 16464 41564 16516
rect 41052 16396 41104 16448
rect 41328 16396 41380 16448
rect 44088 16464 44140 16516
rect 48412 16736 48464 16788
rect 50160 16779 50212 16788
rect 50160 16745 50169 16779
rect 50169 16745 50203 16779
rect 50203 16745 50212 16779
rect 50160 16736 50212 16745
rect 52460 16736 52512 16788
rect 54300 16779 54352 16788
rect 47768 16600 47820 16652
rect 51356 16668 51408 16720
rect 49148 16600 49200 16652
rect 50620 16643 50672 16652
rect 50620 16609 50629 16643
rect 50629 16609 50663 16643
rect 50663 16609 50672 16643
rect 50620 16600 50672 16609
rect 51448 16643 51500 16652
rect 51448 16609 51457 16643
rect 51457 16609 51491 16643
rect 51491 16609 51500 16643
rect 51448 16600 51500 16609
rect 52828 16668 52880 16720
rect 53380 16668 53432 16720
rect 54300 16745 54309 16779
rect 54309 16745 54343 16779
rect 54343 16745 54352 16779
rect 54300 16736 54352 16745
rect 48320 16575 48372 16584
rect 48320 16541 48329 16575
rect 48329 16541 48363 16575
rect 48363 16541 48372 16575
rect 48320 16532 48372 16541
rect 49056 16532 49108 16584
rect 52000 16532 52052 16584
rect 52460 16464 52512 16516
rect 43904 16439 43956 16448
rect 43904 16405 43913 16439
rect 43913 16405 43947 16439
rect 43947 16405 43956 16439
rect 43904 16396 43956 16405
rect 45836 16396 45888 16448
rect 48136 16439 48188 16448
rect 48136 16405 48145 16439
rect 48145 16405 48179 16439
rect 48179 16405 48188 16439
rect 48136 16396 48188 16405
rect 48228 16396 48280 16448
rect 49240 16396 49292 16448
rect 52736 16439 52788 16448
rect 52736 16405 52745 16439
rect 52745 16405 52779 16439
rect 52779 16405 52788 16439
rect 52736 16396 52788 16405
rect 52828 16396 52880 16448
rect 53288 16532 53340 16584
rect 54392 16600 54444 16652
rect 55404 16643 55456 16652
rect 55404 16609 55413 16643
rect 55413 16609 55447 16643
rect 55447 16609 55456 16643
rect 55404 16600 55456 16609
rect 56324 16600 56376 16652
rect 56692 16643 56744 16652
rect 56692 16609 56701 16643
rect 56701 16609 56735 16643
rect 56735 16609 56744 16643
rect 56692 16600 56744 16609
rect 53932 16575 53984 16584
rect 53932 16541 53941 16575
rect 53941 16541 53975 16575
rect 53975 16541 53984 16575
rect 53932 16532 53984 16541
rect 55220 16532 55272 16584
rect 55496 16575 55548 16584
rect 55496 16541 55505 16575
rect 55505 16541 55539 16575
rect 55539 16541 55548 16575
rect 55496 16532 55548 16541
rect 53196 16464 53248 16516
rect 57428 16464 57480 16516
rect 54116 16396 54168 16448
rect 56600 16396 56652 16448
rect 56784 16396 56836 16448
rect 15398 16294 15450 16346
rect 15462 16294 15514 16346
rect 15526 16294 15578 16346
rect 15590 16294 15642 16346
rect 15654 16294 15706 16346
rect 29846 16294 29898 16346
rect 29910 16294 29962 16346
rect 29974 16294 30026 16346
rect 30038 16294 30090 16346
rect 30102 16294 30154 16346
rect 44294 16294 44346 16346
rect 44358 16294 44410 16346
rect 44422 16294 44474 16346
rect 44486 16294 44538 16346
rect 44550 16294 44602 16346
rect 3424 16235 3476 16244
rect 3424 16201 3433 16235
rect 3433 16201 3467 16235
rect 3467 16201 3476 16235
rect 3424 16192 3476 16201
rect 9864 16192 9916 16244
rect 14280 16192 14332 16244
rect 18972 16192 19024 16244
rect 3332 16124 3384 16176
rect 4068 16056 4120 16108
rect 6736 16124 6788 16176
rect 9956 16124 10008 16176
rect 12256 16167 12308 16176
rect 12256 16133 12265 16167
rect 12265 16133 12299 16167
rect 12299 16133 12308 16167
rect 12256 16124 12308 16133
rect 12716 16124 12768 16176
rect 15752 16124 15804 16176
rect 19708 16167 19760 16176
rect 19708 16133 19717 16167
rect 19717 16133 19751 16167
rect 19751 16133 19760 16167
rect 19708 16124 19760 16133
rect 20168 16124 20220 16176
rect 5264 16056 5316 16108
rect 7196 16056 7248 16108
rect 14372 16099 14424 16108
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 14372 16065 14381 16099
rect 14381 16065 14415 16099
rect 14415 16065 14424 16099
rect 14372 16056 14424 16065
rect 22284 16056 22336 16108
rect 23112 16192 23164 16244
rect 23204 16167 23256 16176
rect 23204 16133 23213 16167
rect 23213 16133 23247 16167
rect 23247 16133 23256 16167
rect 23204 16124 23256 16133
rect 24492 16124 24544 16176
rect 10600 15988 10652 16040
rect 10692 15988 10744 16040
rect 11980 16031 12032 16040
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 12992 15988 13044 16040
rect 16304 15988 16356 16040
rect 17224 16031 17276 16040
rect 17224 15997 17233 16031
rect 17233 15997 17267 16031
rect 17267 15997 17276 16031
rect 17224 15988 17276 15997
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 19432 16031 19484 16040
rect 5816 15963 5868 15972
rect 5816 15929 5825 15963
rect 5825 15929 5859 15963
rect 5859 15929 5868 15963
rect 5816 15920 5868 15929
rect 6460 15963 6512 15972
rect 6460 15929 6469 15963
rect 6469 15929 6503 15963
rect 6503 15929 6512 15963
rect 6460 15920 6512 15929
rect 6736 15920 6788 15972
rect 14740 15920 14792 15972
rect 19432 15997 19441 16031
rect 19441 15997 19475 16031
rect 19475 15997 19484 16031
rect 19432 15988 19484 15997
rect 20260 15988 20312 16040
rect 29736 16192 29788 16244
rect 31760 16192 31812 16244
rect 24676 16124 24728 16176
rect 28080 16124 28132 16176
rect 37648 16192 37700 16244
rect 26608 16056 26660 16108
rect 27620 16099 27672 16108
rect 27620 16065 27629 16099
rect 27629 16065 27663 16099
rect 27663 16065 27672 16099
rect 27620 16056 27672 16065
rect 34060 16124 34112 16176
rect 35256 16124 35308 16176
rect 39396 16192 39448 16244
rect 41696 16192 41748 16244
rect 27712 16031 27764 16040
rect 27712 15997 27721 16031
rect 27721 15997 27755 16031
rect 27755 15997 27764 16031
rect 27712 15988 27764 15997
rect 7932 15852 7984 15904
rect 8852 15852 8904 15904
rect 15292 15852 15344 15904
rect 16120 15852 16172 15904
rect 20996 15852 21048 15904
rect 21088 15852 21140 15904
rect 27344 15920 27396 15972
rect 27528 15920 27580 15972
rect 30932 16056 30984 16108
rect 29276 15988 29328 16040
rect 30564 15988 30616 16040
rect 32128 16031 32180 16040
rect 32128 15997 32137 16031
rect 32137 15997 32171 16031
rect 32171 15997 32180 16031
rect 32128 15988 32180 15997
rect 32404 16031 32456 16040
rect 32404 15997 32413 16031
rect 32413 15997 32447 16031
rect 32447 15997 32456 16031
rect 32404 15988 32456 15997
rect 33140 15988 33192 16040
rect 36268 16056 36320 16108
rect 42064 16124 42116 16176
rect 38568 16099 38620 16108
rect 35808 15988 35860 16040
rect 36176 15988 36228 16040
rect 38568 16065 38577 16099
rect 38577 16065 38611 16099
rect 38611 16065 38620 16099
rect 38568 16056 38620 16065
rect 39028 16099 39080 16108
rect 39028 16065 39037 16099
rect 39037 16065 39071 16099
rect 39071 16065 39080 16099
rect 39028 16056 39080 16065
rect 39672 16099 39724 16108
rect 39672 16065 39681 16099
rect 39681 16065 39715 16099
rect 39715 16065 39724 16099
rect 39672 16056 39724 16065
rect 41052 16099 41104 16108
rect 41052 16065 41061 16099
rect 41061 16065 41095 16099
rect 41095 16065 41104 16099
rect 41052 16056 41104 16065
rect 45652 16192 45704 16244
rect 46848 16192 46900 16244
rect 48136 16192 48188 16244
rect 50068 16192 50120 16244
rect 52460 16192 52512 16244
rect 54208 16192 54260 16244
rect 55404 16192 55456 16244
rect 45192 16124 45244 16176
rect 45560 16167 45612 16176
rect 45560 16133 45569 16167
rect 45569 16133 45603 16167
rect 45603 16133 45612 16167
rect 45560 16124 45612 16133
rect 45836 16099 45888 16108
rect 45836 16065 45845 16099
rect 45845 16065 45879 16099
rect 45879 16065 45888 16099
rect 45836 16056 45888 16065
rect 46480 16099 46532 16108
rect 46480 16065 46489 16099
rect 46489 16065 46523 16099
rect 46523 16065 46532 16099
rect 46480 16056 46532 16065
rect 48964 16124 49016 16176
rect 41236 15988 41288 16040
rect 41880 16031 41932 16040
rect 41880 15997 41889 16031
rect 41889 15997 41923 16031
rect 41923 15997 41932 16031
rect 41880 15988 41932 15997
rect 33876 15920 33928 15972
rect 38844 15920 38896 15972
rect 39028 15920 39080 15972
rect 44180 15988 44232 16040
rect 46756 16031 46808 16040
rect 46756 15997 46765 16031
rect 46765 15997 46799 16031
rect 46799 15997 46808 16031
rect 48136 16056 48188 16108
rect 48320 16056 48372 16108
rect 46756 15988 46808 15997
rect 48044 15988 48096 16040
rect 49332 16056 49384 16108
rect 51356 16056 51408 16108
rect 52736 16099 52788 16108
rect 52736 16065 52745 16099
rect 52745 16065 52779 16099
rect 52779 16065 52788 16099
rect 52736 16056 52788 16065
rect 53380 16124 53432 16176
rect 53564 16124 53616 16176
rect 54116 16056 54168 16108
rect 54760 16099 54812 16108
rect 54760 16065 54769 16099
rect 54769 16065 54803 16099
rect 54803 16065 54812 16099
rect 54760 16056 54812 16065
rect 54944 16099 54996 16108
rect 54944 16065 54953 16099
rect 54953 16065 54987 16099
rect 54987 16065 54996 16099
rect 54944 16056 54996 16065
rect 46020 15920 46072 15972
rect 48228 15920 48280 15972
rect 52552 15988 52604 16040
rect 55036 15988 55088 16040
rect 55772 16099 55824 16108
rect 55772 16065 55781 16099
rect 55781 16065 55815 16099
rect 55815 16065 55824 16099
rect 55772 16056 55824 16065
rect 56416 16056 56468 16108
rect 57152 16099 57204 16108
rect 57152 16065 57161 16099
rect 57161 16065 57195 16099
rect 57195 16065 57204 16099
rect 57152 16056 57204 16065
rect 57060 16031 57112 16040
rect 57060 15997 57069 16031
rect 57069 15997 57103 16031
rect 57103 15997 57112 16031
rect 57060 15988 57112 15997
rect 24400 15852 24452 15904
rect 25412 15852 25464 15904
rect 30380 15852 30432 15904
rect 34888 15852 34940 15904
rect 38568 15895 38620 15904
rect 38568 15861 38577 15895
rect 38577 15861 38611 15895
rect 38611 15861 38620 15895
rect 38568 15852 38620 15861
rect 44732 15852 44784 15904
rect 45008 15852 45060 15904
rect 45560 15852 45612 15904
rect 48320 15852 48372 15904
rect 53196 15920 53248 15972
rect 56692 15920 56744 15972
rect 49700 15895 49752 15904
rect 49700 15861 49709 15895
rect 49709 15861 49743 15895
rect 49743 15861 49752 15895
rect 49700 15852 49752 15861
rect 51264 15852 51316 15904
rect 53748 15852 53800 15904
rect 8174 15750 8226 15802
rect 8238 15750 8290 15802
rect 8302 15750 8354 15802
rect 8366 15750 8418 15802
rect 8430 15750 8482 15802
rect 22622 15750 22674 15802
rect 22686 15750 22738 15802
rect 22750 15750 22802 15802
rect 22814 15750 22866 15802
rect 22878 15750 22930 15802
rect 37070 15750 37122 15802
rect 37134 15750 37186 15802
rect 37198 15750 37250 15802
rect 37262 15750 37314 15802
rect 37326 15750 37378 15802
rect 51518 15750 51570 15802
rect 51582 15750 51634 15802
rect 51646 15750 51698 15802
rect 51710 15750 51762 15802
rect 51774 15750 51826 15802
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 10600 15648 10652 15700
rect 10968 15648 11020 15700
rect 16488 15648 16540 15700
rect 18604 15691 18656 15700
rect 18604 15657 18613 15691
rect 18613 15657 18647 15691
rect 18647 15657 18656 15691
rect 18604 15648 18656 15657
rect 20628 15648 20680 15700
rect 23848 15691 23900 15700
rect 23848 15657 23857 15691
rect 23857 15657 23891 15691
rect 23891 15657 23900 15691
rect 23848 15648 23900 15657
rect 24492 15691 24544 15700
rect 24492 15657 24501 15691
rect 24501 15657 24535 15691
rect 24535 15657 24544 15691
rect 24492 15648 24544 15657
rect 5632 15580 5684 15632
rect 6184 15512 6236 15564
rect 8300 15555 8352 15564
rect 8300 15521 8309 15555
rect 8309 15521 8343 15555
rect 8343 15521 8352 15555
rect 8300 15512 8352 15521
rect 8760 15512 8812 15564
rect 5448 15487 5500 15496
rect 5448 15453 5457 15487
rect 5457 15453 5491 15487
rect 5491 15453 5500 15487
rect 5448 15444 5500 15453
rect 6092 15444 6144 15496
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 6736 15487 6788 15496
rect 6736 15453 6745 15487
rect 6745 15453 6779 15487
rect 6779 15453 6788 15487
rect 6736 15444 6788 15453
rect 9128 15444 9180 15496
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 11060 15580 11112 15632
rect 9496 15512 9548 15564
rect 12992 15512 13044 15564
rect 19432 15580 19484 15632
rect 26240 15648 26292 15700
rect 32404 15648 32456 15700
rect 36360 15648 36412 15700
rect 36544 15648 36596 15700
rect 41880 15648 41932 15700
rect 9220 15444 9272 15453
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 10876 15444 10928 15496
rect 12072 15444 12124 15496
rect 18788 15512 18840 15564
rect 20076 15555 20128 15564
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 32036 15580 32088 15632
rect 32220 15580 32272 15632
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 15200 15444 15252 15496
rect 19524 15444 19576 15496
rect 19800 15487 19852 15496
rect 19800 15453 19809 15487
rect 19809 15453 19843 15487
rect 19843 15453 19852 15487
rect 19800 15444 19852 15453
rect 24308 15512 24360 15564
rect 8668 15376 8720 15428
rect 6000 15351 6052 15360
rect 6000 15317 6009 15351
rect 6009 15317 6043 15351
rect 6043 15317 6052 15351
rect 6000 15308 6052 15317
rect 7564 15351 7616 15360
rect 7564 15317 7573 15351
rect 7573 15317 7607 15351
rect 7607 15317 7616 15351
rect 7564 15308 7616 15317
rect 13912 15376 13964 15428
rect 16672 15419 16724 15428
rect 16672 15385 16681 15419
rect 16681 15385 16715 15419
rect 16715 15385 16724 15419
rect 16672 15376 16724 15385
rect 23020 15487 23072 15496
rect 23020 15453 23029 15487
rect 23029 15453 23063 15487
rect 23063 15453 23072 15487
rect 23020 15444 23072 15453
rect 24032 15444 24084 15496
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 22284 15376 22336 15428
rect 23480 15376 23532 15428
rect 13820 15308 13872 15360
rect 24676 15308 24728 15360
rect 27528 15444 27580 15496
rect 29460 15512 29512 15564
rect 33600 15512 33652 15564
rect 36084 15580 36136 15632
rect 29552 15487 29604 15496
rect 29552 15453 29561 15487
rect 29561 15453 29595 15487
rect 29595 15453 29604 15487
rect 29552 15444 29604 15453
rect 33140 15487 33192 15496
rect 33140 15453 33149 15487
rect 33149 15453 33183 15487
rect 33183 15453 33192 15487
rect 33140 15444 33192 15453
rect 33968 15487 34020 15496
rect 33968 15453 33977 15487
rect 33977 15453 34011 15487
rect 34011 15453 34020 15487
rect 38660 15512 38712 15564
rect 39672 15580 39724 15632
rect 38844 15512 38896 15564
rect 39948 15555 40000 15564
rect 39948 15521 39957 15555
rect 39957 15521 39991 15555
rect 39991 15521 40000 15555
rect 39948 15512 40000 15521
rect 47676 15648 47728 15700
rect 49700 15648 49752 15700
rect 51172 15691 51224 15700
rect 51172 15657 51181 15691
rect 51181 15657 51215 15691
rect 51215 15657 51224 15691
rect 51172 15648 51224 15657
rect 53380 15648 53432 15700
rect 54760 15648 54812 15700
rect 55496 15648 55548 15700
rect 44640 15580 44692 15632
rect 48136 15580 48188 15632
rect 45928 15555 45980 15564
rect 33968 15444 34020 15453
rect 37648 15487 37700 15496
rect 37648 15453 37657 15487
rect 37657 15453 37691 15487
rect 37691 15453 37700 15487
rect 37648 15444 37700 15453
rect 38936 15444 38988 15496
rect 40868 15487 40920 15496
rect 40868 15453 40877 15487
rect 40877 15453 40911 15487
rect 40911 15453 40920 15487
rect 40868 15444 40920 15453
rect 44088 15487 44140 15496
rect 44088 15453 44097 15487
rect 44097 15453 44131 15487
rect 44131 15453 44140 15487
rect 44088 15444 44140 15453
rect 27988 15376 28040 15428
rect 29092 15376 29144 15428
rect 31392 15419 31444 15428
rect 31392 15385 31401 15419
rect 31401 15385 31435 15419
rect 31435 15385 31444 15419
rect 31392 15376 31444 15385
rect 31576 15376 31628 15428
rect 32404 15376 32456 15428
rect 35256 15376 35308 15428
rect 26608 15308 26660 15360
rect 28816 15308 28868 15360
rect 32220 15308 32272 15360
rect 38384 15376 38436 15428
rect 41880 15419 41932 15428
rect 41880 15385 41889 15419
rect 41889 15385 41923 15419
rect 41923 15385 41932 15419
rect 41880 15376 41932 15385
rect 45928 15521 45937 15555
rect 45937 15521 45971 15555
rect 45971 15521 45980 15555
rect 45928 15512 45980 15521
rect 46020 15512 46072 15564
rect 48228 15555 48280 15564
rect 45008 15487 45060 15496
rect 45008 15453 45017 15487
rect 45017 15453 45051 15487
rect 45051 15453 45060 15487
rect 45008 15444 45060 15453
rect 48228 15521 48237 15555
rect 48237 15521 48271 15555
rect 48271 15521 48280 15555
rect 48228 15512 48280 15521
rect 49240 15512 49292 15564
rect 36544 15308 36596 15360
rect 38752 15308 38804 15360
rect 46112 15376 46164 15428
rect 46940 15376 46992 15428
rect 47492 15419 47544 15428
rect 47492 15385 47501 15419
rect 47501 15385 47535 15419
rect 47535 15385 47544 15419
rect 47492 15376 47544 15385
rect 49792 15444 49844 15496
rect 51080 15487 51132 15496
rect 51080 15453 51089 15487
rect 51089 15453 51123 15487
rect 51123 15453 51132 15487
rect 51264 15487 51316 15496
rect 51080 15444 51132 15453
rect 51264 15453 51273 15487
rect 51273 15453 51307 15487
rect 51307 15453 51316 15487
rect 51264 15444 51316 15453
rect 54944 15580 54996 15632
rect 52828 15512 52880 15564
rect 56324 15555 56376 15564
rect 56324 15521 56333 15555
rect 56333 15521 56367 15555
rect 56367 15521 56376 15555
rect 56324 15512 56376 15521
rect 56600 15555 56652 15564
rect 56600 15521 56609 15555
rect 56609 15521 56643 15555
rect 56643 15521 56652 15555
rect 56600 15512 56652 15521
rect 52184 15487 52236 15496
rect 52184 15453 52193 15487
rect 52193 15453 52227 15487
rect 52227 15453 52236 15487
rect 52184 15444 52236 15453
rect 49332 15419 49384 15428
rect 44640 15308 44692 15360
rect 44824 15308 44876 15360
rect 45928 15308 45980 15360
rect 47308 15308 47360 15360
rect 48136 15308 48188 15360
rect 48688 15351 48740 15360
rect 48688 15317 48697 15351
rect 48697 15317 48731 15351
rect 48731 15317 48740 15351
rect 48688 15308 48740 15317
rect 49332 15385 49341 15419
rect 49341 15385 49375 15419
rect 49375 15385 49384 15419
rect 49332 15376 49384 15385
rect 50712 15376 50764 15428
rect 53840 15444 53892 15496
rect 52736 15376 52788 15428
rect 53196 15419 53248 15428
rect 53196 15385 53205 15419
rect 53205 15385 53239 15419
rect 53239 15385 53248 15419
rect 53196 15376 53248 15385
rect 53564 15376 53616 15428
rect 54116 15444 54168 15496
rect 54208 15487 54260 15496
rect 54208 15453 54217 15487
rect 54217 15453 54251 15487
rect 54251 15453 54260 15487
rect 54208 15444 54260 15453
rect 55772 15444 55824 15496
rect 57336 15376 57388 15428
rect 49240 15308 49292 15360
rect 49976 15308 50028 15360
rect 51908 15308 51960 15360
rect 52828 15351 52880 15360
rect 52828 15317 52837 15351
rect 52837 15317 52871 15351
rect 52871 15317 52880 15351
rect 52828 15308 52880 15317
rect 53656 15308 53708 15360
rect 15398 15206 15450 15258
rect 15462 15206 15514 15258
rect 15526 15206 15578 15258
rect 15590 15206 15642 15258
rect 15654 15206 15706 15258
rect 29846 15206 29898 15258
rect 29910 15206 29962 15258
rect 29974 15206 30026 15258
rect 30038 15206 30090 15258
rect 30102 15206 30154 15258
rect 44294 15206 44346 15258
rect 44358 15206 44410 15258
rect 44422 15206 44474 15258
rect 44486 15206 44538 15258
rect 44550 15206 44602 15258
rect 5356 15104 5408 15156
rect 6828 15104 6880 15156
rect 10876 15104 10928 15156
rect 15200 15104 15252 15156
rect 12532 15036 12584 15088
rect 15292 15036 15344 15088
rect 5264 14968 5316 15020
rect 6368 14968 6420 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 7932 15011 7984 15020
rect 7932 14977 7941 15011
rect 7941 14977 7975 15011
rect 7975 14977 7984 15011
rect 7932 14968 7984 14977
rect 19432 15104 19484 15156
rect 20168 15104 20220 15156
rect 19248 15036 19300 15088
rect 21088 15104 21140 15156
rect 21364 15104 21416 15156
rect 20720 15036 20772 15088
rect 21824 15079 21876 15088
rect 21824 15045 21833 15079
rect 21833 15045 21867 15079
rect 21867 15045 21876 15079
rect 21824 15036 21876 15045
rect 16764 15011 16816 15020
rect 10600 14900 10652 14952
rect 10692 14900 10744 14952
rect 6552 14832 6604 14884
rect 7840 14764 7892 14816
rect 8024 14807 8076 14816
rect 8024 14773 8033 14807
rect 8033 14773 8067 14807
rect 8067 14773 8076 14807
rect 8024 14764 8076 14773
rect 9680 14764 9732 14816
rect 16764 14977 16773 15011
rect 16773 14977 16807 15011
rect 16807 14977 16816 15011
rect 16764 14968 16816 14977
rect 20812 14968 20864 15020
rect 21088 14968 21140 15020
rect 22192 15036 22244 15088
rect 24676 15079 24728 15088
rect 24676 15045 24685 15079
rect 24685 15045 24719 15079
rect 24719 15045 24728 15079
rect 24676 15036 24728 15045
rect 26976 15104 27028 15156
rect 30472 15104 30524 15156
rect 32128 15104 32180 15156
rect 35164 15104 35216 15156
rect 35440 15104 35492 15156
rect 35992 15147 36044 15156
rect 35992 15113 36001 15147
rect 36001 15113 36035 15147
rect 36035 15113 36044 15147
rect 35992 15104 36044 15113
rect 24032 15011 24084 15020
rect 24032 14977 24041 15011
rect 24041 14977 24075 15011
rect 24075 14977 24084 15011
rect 24032 14968 24084 14977
rect 27804 15036 27856 15088
rect 28632 15036 28684 15088
rect 30564 15079 30616 15088
rect 30564 15045 30573 15079
rect 30573 15045 30607 15079
rect 30607 15045 30616 15079
rect 30564 15036 30616 15045
rect 35256 15036 35308 15088
rect 39948 15104 40000 15156
rect 38752 15079 38804 15088
rect 38752 15045 38761 15079
rect 38761 15045 38795 15079
rect 38795 15045 38804 15079
rect 38752 15036 38804 15045
rect 27620 14968 27672 15020
rect 32312 15011 32364 15020
rect 32312 14977 32321 15011
rect 32321 14977 32355 15011
rect 32355 14977 32364 15011
rect 32312 14968 32364 14977
rect 33600 15011 33652 15020
rect 33600 14977 33609 15011
rect 33609 14977 33643 15011
rect 33643 14977 33652 15011
rect 33600 14968 33652 14977
rect 36452 14968 36504 15020
rect 12532 14900 12584 14952
rect 17500 14943 17552 14952
rect 12256 14764 12308 14816
rect 14004 14764 14056 14816
rect 17500 14909 17509 14943
rect 17509 14909 17543 14943
rect 17543 14909 17552 14943
rect 17500 14900 17552 14909
rect 18972 14943 19024 14952
rect 18972 14909 18981 14943
rect 18981 14909 19015 14943
rect 19015 14909 19024 14943
rect 18972 14900 19024 14909
rect 19708 14900 19760 14952
rect 21640 14900 21692 14952
rect 21916 14900 21968 14952
rect 19524 14832 19576 14884
rect 23572 14900 23624 14952
rect 29092 14900 29144 14952
rect 33048 14900 33100 14952
rect 33232 14900 33284 14952
rect 26976 14832 27028 14884
rect 19892 14764 19944 14816
rect 24216 14807 24268 14816
rect 24216 14773 24225 14807
rect 24225 14773 24259 14807
rect 24259 14773 24268 14807
rect 24216 14764 24268 14773
rect 25964 14807 26016 14816
rect 25964 14773 25973 14807
rect 25973 14773 26007 14807
rect 26007 14773 26016 14807
rect 25964 14764 26016 14773
rect 28080 14807 28132 14816
rect 28080 14773 28089 14807
rect 28089 14773 28123 14807
rect 28123 14773 28132 14807
rect 28080 14764 28132 14773
rect 32220 14807 32272 14816
rect 32220 14773 32229 14807
rect 32229 14773 32263 14807
rect 32263 14773 32272 14807
rect 32220 14764 32272 14773
rect 36636 14807 36688 14816
rect 36636 14773 36645 14807
rect 36645 14773 36679 14807
rect 36679 14773 36688 14807
rect 36636 14764 36688 14773
rect 39028 15011 39080 15020
rect 39028 14977 39037 15011
rect 39037 14977 39071 15011
rect 39071 14977 39080 15011
rect 39028 14968 39080 14977
rect 40132 14968 40184 15020
rect 40684 15104 40736 15156
rect 45008 15104 45060 15156
rect 45468 15104 45520 15156
rect 50712 15147 50764 15156
rect 40500 14900 40552 14952
rect 41420 15036 41472 15088
rect 41880 15036 41932 15088
rect 41144 14968 41196 15020
rect 41788 14968 41840 15020
rect 44732 15036 44784 15088
rect 46848 15036 46900 15088
rect 47492 14968 47544 15020
rect 41420 14900 41472 14952
rect 42616 14900 42668 14952
rect 42892 14900 42944 14952
rect 44824 14943 44876 14952
rect 44824 14909 44833 14943
rect 44833 14909 44867 14943
rect 44867 14909 44876 14943
rect 44824 14900 44876 14909
rect 45100 14943 45152 14952
rect 45100 14909 45109 14943
rect 45109 14909 45143 14943
rect 45143 14909 45152 14943
rect 45100 14900 45152 14909
rect 45836 14900 45888 14952
rect 50712 15113 50721 15147
rect 50721 15113 50755 15147
rect 50755 15113 50764 15147
rect 50712 15104 50764 15113
rect 52184 15104 52236 15156
rect 48688 15036 48740 15088
rect 50252 15036 50304 15088
rect 52828 15036 52880 15088
rect 51356 15011 51408 15020
rect 51356 14977 51365 15011
rect 51365 14977 51399 15011
rect 51399 14977 51408 15011
rect 51356 14968 51408 14977
rect 44640 14832 44692 14884
rect 48228 14900 48280 14952
rect 49792 14900 49844 14952
rect 51448 14943 51500 14952
rect 51448 14909 51457 14943
rect 51457 14909 51491 14943
rect 51491 14909 51500 14943
rect 51448 14900 51500 14909
rect 53104 14968 53156 15020
rect 53288 14968 53340 15020
rect 56048 15036 56100 15088
rect 38292 14764 38344 14816
rect 42984 14764 43036 14816
rect 44916 14764 44968 14816
rect 48872 14832 48924 14884
rect 48044 14807 48096 14816
rect 48044 14773 48053 14807
rect 48053 14773 48087 14807
rect 48087 14773 48096 14807
rect 48044 14764 48096 14773
rect 49700 14764 49752 14816
rect 51264 14764 51316 14816
rect 53472 14900 53524 14952
rect 53748 14900 53800 14952
rect 56876 14943 56928 14952
rect 56876 14909 56885 14943
rect 56885 14909 56919 14943
rect 56919 14909 56928 14943
rect 56876 14900 56928 14909
rect 53380 14764 53432 14816
rect 57152 14764 57204 14816
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 8302 14662 8354 14714
rect 8366 14662 8418 14714
rect 8430 14662 8482 14714
rect 22622 14662 22674 14714
rect 22686 14662 22738 14714
rect 22750 14662 22802 14714
rect 22814 14662 22866 14714
rect 22878 14662 22930 14714
rect 37070 14662 37122 14714
rect 37134 14662 37186 14714
rect 37198 14662 37250 14714
rect 37262 14662 37314 14714
rect 37326 14662 37378 14714
rect 51518 14662 51570 14714
rect 51582 14662 51634 14714
rect 51646 14662 51698 14714
rect 51710 14662 51762 14714
rect 51774 14662 51826 14714
rect 5264 14560 5316 14612
rect 6644 14560 6696 14612
rect 8852 14560 8904 14612
rect 9956 14560 10008 14612
rect 10600 14560 10652 14612
rect 13912 14560 13964 14612
rect 14740 14560 14792 14612
rect 19248 14560 19300 14612
rect 19800 14560 19852 14612
rect 19892 14560 19944 14612
rect 23572 14560 23624 14612
rect 8300 14535 8352 14544
rect 8300 14501 8309 14535
rect 8309 14501 8343 14535
rect 8343 14501 8352 14535
rect 8300 14492 8352 14501
rect 8944 14492 8996 14544
rect 10876 14492 10928 14544
rect 14372 14492 14424 14544
rect 19340 14492 19392 14544
rect 5908 14424 5960 14476
rect 7932 14424 7984 14476
rect 8668 14356 8720 14408
rect 9680 14356 9732 14408
rect 9864 14424 9916 14476
rect 15752 14424 15804 14476
rect 7748 14220 7800 14272
rect 10600 14220 10652 14272
rect 12808 14356 12860 14408
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 16028 14399 16080 14408
rect 16028 14365 16037 14399
rect 16037 14365 16071 14399
rect 16071 14365 16080 14399
rect 18512 14424 18564 14476
rect 16488 14399 16540 14408
rect 16028 14356 16080 14365
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 17132 14356 17184 14408
rect 19524 14399 19576 14408
rect 12440 14288 12492 14340
rect 13820 14288 13872 14340
rect 17316 14288 17368 14340
rect 19524 14365 19533 14399
rect 19533 14365 19567 14399
rect 19567 14365 19576 14399
rect 19524 14356 19576 14365
rect 21180 14467 21232 14476
rect 21180 14433 21189 14467
rect 21189 14433 21223 14467
rect 21223 14433 21232 14467
rect 21180 14424 21232 14433
rect 23940 14424 23992 14476
rect 24768 14560 24820 14612
rect 27344 14560 27396 14612
rect 29000 14603 29052 14612
rect 27620 14492 27672 14544
rect 29000 14569 29009 14603
rect 29009 14569 29043 14603
rect 29043 14569 29052 14603
rect 29000 14560 29052 14569
rect 33968 14560 34020 14612
rect 28080 14424 28132 14476
rect 30472 14424 30524 14476
rect 32312 14492 32364 14544
rect 37096 14560 37148 14612
rect 36636 14467 36688 14476
rect 36636 14433 36645 14467
rect 36645 14433 36679 14467
rect 36679 14433 36688 14467
rect 36636 14424 36688 14433
rect 38660 14424 38712 14476
rect 45100 14560 45152 14612
rect 46112 14603 46164 14612
rect 46112 14569 46121 14603
rect 46121 14569 46155 14603
rect 46155 14569 46164 14603
rect 46112 14560 46164 14569
rect 48780 14560 48832 14612
rect 48872 14560 48924 14612
rect 52920 14560 52972 14612
rect 42524 14492 42576 14544
rect 43996 14492 44048 14544
rect 44180 14492 44232 14544
rect 45376 14535 45428 14544
rect 45376 14501 45385 14535
rect 45385 14501 45419 14535
rect 45419 14501 45428 14535
rect 45376 14492 45428 14501
rect 45836 14492 45888 14544
rect 20812 14356 20864 14408
rect 21272 14356 21324 14408
rect 22008 14356 22060 14408
rect 23480 14356 23532 14408
rect 26792 14399 26844 14408
rect 26792 14365 26801 14399
rect 26801 14365 26835 14399
rect 26835 14365 26844 14399
rect 26792 14356 26844 14365
rect 27436 14399 27488 14408
rect 27436 14365 27445 14399
rect 27445 14365 27479 14399
rect 27479 14365 27488 14399
rect 27436 14356 27488 14365
rect 27620 14399 27672 14408
rect 27620 14365 27629 14399
rect 27629 14365 27663 14399
rect 27663 14365 27672 14399
rect 27620 14356 27672 14365
rect 29736 14356 29788 14408
rect 20168 14288 20220 14340
rect 20260 14288 20312 14340
rect 21916 14288 21968 14340
rect 22376 14331 22428 14340
rect 22376 14297 22385 14331
rect 22385 14297 22419 14331
rect 22419 14297 22428 14331
rect 22376 14288 22428 14297
rect 25412 14288 25464 14340
rect 32220 14288 32272 14340
rect 36544 14288 36596 14340
rect 12348 14220 12400 14272
rect 14372 14220 14424 14272
rect 18512 14220 18564 14272
rect 21364 14220 21416 14272
rect 22192 14220 22244 14272
rect 23020 14220 23072 14272
rect 26700 14263 26752 14272
rect 26700 14229 26709 14263
rect 26709 14229 26743 14263
rect 26743 14229 26752 14263
rect 26700 14220 26752 14229
rect 28448 14263 28500 14272
rect 28448 14229 28457 14263
rect 28457 14229 28491 14263
rect 28491 14229 28500 14263
rect 28448 14220 28500 14229
rect 32588 14220 32640 14272
rect 37648 14356 37700 14408
rect 38292 14399 38344 14408
rect 38292 14365 38301 14399
rect 38301 14365 38335 14399
rect 38335 14365 38344 14399
rect 38292 14356 38344 14365
rect 40592 14356 40644 14408
rect 40684 14356 40736 14408
rect 41144 14356 41196 14408
rect 41420 14356 41472 14408
rect 39304 14288 39356 14340
rect 41696 14356 41748 14408
rect 44916 14424 44968 14476
rect 46204 14467 46256 14476
rect 46204 14433 46213 14467
rect 46213 14433 46247 14467
rect 46247 14433 46256 14467
rect 46204 14424 46256 14433
rect 46296 14424 46348 14476
rect 48964 14492 49016 14544
rect 42892 14399 42944 14408
rect 41788 14288 41840 14340
rect 42524 14288 42576 14340
rect 42892 14365 42901 14399
rect 42901 14365 42935 14399
rect 42935 14365 42944 14399
rect 42892 14356 42944 14365
rect 43536 14399 43588 14408
rect 43536 14365 43545 14399
rect 43545 14365 43579 14399
rect 43579 14365 43588 14399
rect 43536 14356 43588 14365
rect 44640 14356 44692 14408
rect 45560 14356 45612 14408
rect 46664 14356 46716 14408
rect 46848 14399 46900 14408
rect 46848 14365 46857 14399
rect 46857 14365 46891 14399
rect 46891 14365 46900 14399
rect 46848 14356 46900 14365
rect 50896 14424 50948 14476
rect 51908 14424 51960 14476
rect 52368 14492 52420 14544
rect 48320 14399 48372 14408
rect 48320 14365 48329 14399
rect 48329 14365 48363 14399
rect 48363 14365 48372 14399
rect 48964 14399 49016 14408
rect 48320 14356 48372 14365
rect 48964 14365 48973 14399
rect 48973 14365 49007 14399
rect 49007 14365 49016 14399
rect 48964 14356 49016 14365
rect 49148 14399 49200 14408
rect 49148 14365 49157 14399
rect 49157 14365 49191 14399
rect 49191 14365 49200 14399
rect 49148 14356 49200 14365
rect 51356 14356 51408 14408
rect 51448 14356 51500 14408
rect 44824 14288 44876 14340
rect 45192 14288 45244 14340
rect 45836 14288 45888 14340
rect 37096 14220 37148 14272
rect 40132 14220 40184 14272
rect 42064 14220 42116 14272
rect 42984 14220 43036 14272
rect 43996 14220 44048 14272
rect 45928 14220 45980 14272
rect 47216 14263 47268 14272
rect 47216 14229 47225 14263
rect 47225 14229 47259 14263
rect 47259 14229 47268 14263
rect 47216 14220 47268 14229
rect 47492 14220 47544 14272
rect 51172 14288 51224 14340
rect 48964 14220 49016 14272
rect 50344 14220 50396 14272
rect 50712 14220 50764 14272
rect 50896 14263 50948 14272
rect 50896 14229 50905 14263
rect 50905 14229 50939 14263
rect 50939 14229 50948 14263
rect 52920 14288 52972 14340
rect 53196 14424 53248 14476
rect 53288 14399 53340 14408
rect 53288 14365 53297 14399
rect 53297 14365 53331 14399
rect 53331 14365 53340 14399
rect 53288 14356 53340 14365
rect 53380 14399 53432 14408
rect 53380 14365 53389 14399
rect 53389 14365 53423 14399
rect 53423 14365 53432 14399
rect 53380 14356 53432 14365
rect 53656 14356 53708 14408
rect 54024 14399 54076 14408
rect 54024 14365 54033 14399
rect 54033 14365 54067 14399
rect 54067 14365 54076 14399
rect 54024 14356 54076 14365
rect 54484 14356 54536 14408
rect 56876 14560 56928 14612
rect 57152 14560 57204 14612
rect 56692 14467 56744 14476
rect 56692 14433 56701 14467
rect 56701 14433 56735 14467
rect 56735 14433 56744 14467
rect 56692 14424 56744 14433
rect 53472 14288 53524 14340
rect 57336 14288 57388 14340
rect 50896 14220 50948 14229
rect 51908 14220 51960 14272
rect 56140 14220 56192 14272
rect 15398 14118 15450 14170
rect 15462 14118 15514 14170
rect 15526 14118 15578 14170
rect 15590 14118 15642 14170
rect 15654 14118 15706 14170
rect 29846 14118 29898 14170
rect 29910 14118 29962 14170
rect 29974 14118 30026 14170
rect 30038 14118 30090 14170
rect 30102 14118 30154 14170
rect 44294 14118 44346 14170
rect 44358 14118 44410 14170
rect 44422 14118 44474 14170
rect 44486 14118 44538 14170
rect 44550 14118 44602 14170
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 11428 14016 11480 14068
rect 8024 13948 8076 14000
rect 10416 13948 10468 14000
rect 11796 14016 11848 14068
rect 12348 14016 12400 14068
rect 6736 13923 6788 13932
rect 6736 13889 6745 13923
rect 6745 13889 6779 13923
rect 6779 13889 6788 13923
rect 6736 13880 6788 13889
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 12348 13880 12400 13932
rect 16028 14016 16080 14068
rect 17132 14016 17184 14068
rect 17316 14059 17368 14068
rect 17316 14025 17325 14059
rect 17325 14025 17359 14059
rect 17359 14025 17368 14059
rect 17316 14016 17368 14025
rect 18512 14059 18564 14068
rect 18512 14025 18521 14059
rect 18521 14025 18555 14059
rect 18555 14025 18564 14059
rect 18512 14016 18564 14025
rect 17960 13948 18012 14000
rect 14004 13880 14056 13932
rect 16580 13880 16632 13932
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 9220 13855 9272 13864
rect 9220 13821 9229 13855
rect 9229 13821 9263 13855
rect 9263 13821 9272 13855
rect 9220 13812 9272 13821
rect 10692 13812 10744 13864
rect 13912 13812 13964 13864
rect 14740 13812 14792 13864
rect 22836 14016 22888 14068
rect 23940 14059 23992 14068
rect 23940 14025 23949 14059
rect 23949 14025 23983 14059
rect 23983 14025 23992 14059
rect 23940 14016 23992 14025
rect 27436 14016 27488 14068
rect 29736 14016 29788 14068
rect 18696 13948 18748 14000
rect 24400 13948 24452 14000
rect 26700 13948 26752 14000
rect 29644 13948 29696 14000
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20260 13880 20312 13889
rect 20996 13880 21048 13932
rect 26240 13880 26292 13932
rect 27804 13923 27856 13932
rect 27804 13889 27813 13923
rect 27813 13889 27847 13923
rect 27847 13889 27856 13923
rect 27804 13880 27856 13889
rect 31024 13880 31076 13932
rect 7840 13744 7892 13796
rect 11428 13744 11480 13796
rect 13544 13744 13596 13796
rect 19984 13812 20036 13864
rect 23204 13812 23256 13864
rect 24124 13812 24176 13864
rect 24768 13812 24820 13864
rect 27068 13855 27120 13864
rect 27068 13821 27077 13855
rect 27077 13821 27111 13855
rect 27111 13821 27120 13855
rect 27068 13812 27120 13821
rect 27528 13812 27580 13864
rect 28080 13855 28132 13864
rect 28080 13821 28089 13855
rect 28089 13821 28123 13855
rect 28123 13821 28132 13855
rect 28080 13812 28132 13821
rect 30748 13812 30800 13864
rect 31208 13923 31260 13932
rect 31208 13889 31217 13923
rect 31217 13889 31251 13923
rect 31251 13889 31260 13923
rect 31208 13880 31260 13889
rect 31300 13812 31352 13864
rect 34244 13948 34296 14000
rect 34888 13948 34940 14000
rect 41696 14016 41748 14068
rect 40684 13948 40736 14000
rect 33600 13880 33652 13932
rect 40040 13923 40092 13932
rect 40040 13889 40049 13923
rect 40049 13889 40083 13923
rect 40083 13889 40092 13923
rect 40040 13880 40092 13889
rect 40960 13923 41012 13932
rect 40960 13889 40969 13923
rect 40969 13889 41003 13923
rect 41003 13889 41012 13923
rect 40960 13880 41012 13889
rect 41696 13923 41748 13932
rect 41696 13889 41705 13923
rect 41705 13889 41739 13923
rect 41739 13889 41748 13923
rect 41696 13880 41748 13889
rect 42524 13948 42576 14000
rect 42708 13923 42760 13932
rect 42708 13889 42717 13923
rect 42717 13889 42751 13923
rect 42751 13889 42760 13923
rect 42708 13880 42760 13889
rect 43996 14016 44048 14068
rect 45468 14016 45520 14068
rect 46296 14016 46348 14068
rect 46664 14059 46716 14068
rect 46664 14025 46673 14059
rect 46673 14025 46707 14059
rect 46707 14025 46716 14059
rect 46664 14016 46716 14025
rect 43444 13948 43496 14000
rect 44824 13991 44876 14000
rect 32680 13855 32732 13864
rect 32680 13821 32689 13855
rect 32689 13821 32723 13855
rect 32723 13821 32732 13855
rect 32680 13812 32732 13821
rect 29092 13744 29144 13796
rect 15844 13676 15896 13728
rect 19616 13676 19668 13728
rect 30196 13676 30248 13728
rect 30380 13719 30432 13728
rect 30380 13685 30389 13719
rect 30389 13685 30423 13719
rect 30423 13685 30432 13719
rect 30380 13676 30432 13685
rect 32404 13744 32456 13796
rect 34244 13812 34296 13864
rect 39304 13812 39356 13864
rect 39396 13855 39448 13864
rect 39396 13821 39405 13855
rect 39405 13821 39439 13855
rect 39439 13821 39448 13855
rect 40684 13855 40736 13864
rect 39396 13812 39448 13821
rect 40684 13821 40693 13855
rect 40693 13821 40727 13855
rect 40727 13821 40736 13855
rect 40684 13812 40736 13821
rect 44824 13957 44833 13991
rect 44833 13957 44867 13991
rect 44867 13957 44876 13991
rect 44824 13948 44876 13957
rect 44916 13948 44968 14000
rect 45100 13991 45152 14000
rect 45100 13957 45109 13991
rect 45109 13957 45143 13991
rect 45143 13957 45152 13991
rect 45100 13948 45152 13957
rect 45192 13923 45244 13932
rect 45192 13889 45201 13923
rect 45201 13889 45235 13923
rect 45235 13889 45244 13923
rect 45192 13880 45244 13889
rect 45836 13923 45888 13932
rect 45836 13889 45845 13923
rect 45845 13889 45879 13923
rect 45879 13889 45888 13923
rect 45836 13880 45888 13889
rect 46020 13880 46072 13932
rect 48044 14016 48096 14068
rect 48228 14016 48280 14068
rect 47216 13948 47268 14000
rect 48136 13948 48188 14000
rect 49240 14016 49292 14068
rect 50620 14059 50672 14068
rect 50620 14025 50629 14059
rect 50629 14025 50663 14059
rect 50663 14025 50672 14059
rect 50620 14016 50672 14025
rect 51264 14016 51316 14068
rect 53840 14059 53892 14068
rect 53840 14025 53849 14059
rect 53849 14025 53883 14059
rect 53883 14025 53892 14059
rect 53840 14016 53892 14025
rect 55588 14016 55640 14068
rect 57244 14059 57296 14068
rect 57244 14025 57253 14059
rect 57253 14025 57287 14059
rect 57287 14025 57296 14059
rect 57244 14016 57296 14025
rect 50896 13948 50948 14000
rect 53472 13948 53524 14000
rect 51172 13880 51224 13932
rect 52184 13880 52236 13932
rect 53196 13923 53248 13932
rect 53196 13889 53205 13923
rect 53205 13889 53239 13923
rect 53239 13889 53248 13923
rect 53196 13880 53248 13889
rect 54024 13923 54076 13932
rect 54024 13889 54033 13923
rect 54033 13889 54067 13923
rect 54067 13889 54076 13923
rect 54024 13880 54076 13889
rect 54208 13880 54260 13932
rect 54484 13923 54536 13932
rect 54484 13889 54493 13923
rect 54493 13889 54527 13923
rect 54527 13889 54536 13923
rect 54484 13880 54536 13889
rect 57980 13880 58032 13932
rect 46204 13812 46256 13864
rect 43536 13744 43588 13796
rect 45928 13787 45980 13796
rect 45928 13753 45937 13787
rect 45937 13753 45971 13787
rect 45971 13753 45980 13787
rect 45928 13744 45980 13753
rect 42156 13676 42208 13728
rect 49976 13812 50028 13864
rect 51356 13855 51408 13864
rect 51356 13821 51365 13855
rect 51365 13821 51399 13855
rect 51399 13821 51408 13855
rect 51356 13812 51408 13821
rect 56140 13855 56192 13864
rect 54208 13744 54260 13796
rect 56140 13821 56149 13855
rect 56149 13821 56183 13855
rect 56183 13821 56192 13855
rect 56140 13812 56192 13821
rect 56048 13744 56100 13796
rect 49148 13676 49200 13728
rect 56692 13676 56744 13728
rect 57888 13719 57940 13728
rect 57888 13685 57897 13719
rect 57897 13685 57931 13719
rect 57931 13685 57940 13719
rect 57888 13676 57940 13685
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 8302 13574 8354 13626
rect 8366 13574 8418 13626
rect 8430 13574 8482 13626
rect 22622 13574 22674 13626
rect 22686 13574 22738 13626
rect 22750 13574 22802 13626
rect 22814 13574 22866 13626
rect 22878 13574 22930 13626
rect 37070 13574 37122 13626
rect 37134 13574 37186 13626
rect 37198 13574 37250 13626
rect 37262 13574 37314 13626
rect 37326 13574 37378 13626
rect 51518 13574 51570 13626
rect 51582 13574 51634 13626
rect 51646 13574 51698 13626
rect 51710 13574 51762 13626
rect 51774 13574 51826 13626
rect 6000 13472 6052 13524
rect 6920 13404 6972 13456
rect 10416 13472 10468 13524
rect 12440 13472 12492 13524
rect 17040 13472 17092 13524
rect 24032 13472 24084 13524
rect 24400 13472 24452 13524
rect 26792 13472 26844 13524
rect 28080 13472 28132 13524
rect 29644 13515 29696 13524
rect 29644 13481 29653 13515
rect 29653 13481 29687 13515
rect 29687 13481 29696 13515
rect 29644 13472 29696 13481
rect 33968 13515 34020 13524
rect 33968 13481 33977 13515
rect 33977 13481 34011 13515
rect 34011 13481 34020 13515
rect 33968 13472 34020 13481
rect 39948 13472 40000 13524
rect 40040 13472 40092 13524
rect 40592 13472 40644 13524
rect 42616 13472 42668 13524
rect 22376 13404 22428 13456
rect 22468 13404 22520 13456
rect 8024 13336 8076 13388
rect 7932 13268 7984 13320
rect 15292 13336 15344 13388
rect 15752 13336 15804 13388
rect 14372 13268 14424 13320
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 24584 13336 24636 13388
rect 30748 13336 30800 13388
rect 16028 13268 16080 13277
rect 13912 13200 13964 13252
rect 16580 13200 16632 13252
rect 8024 13132 8076 13184
rect 13728 13132 13780 13184
rect 14280 13175 14332 13184
rect 14280 13141 14289 13175
rect 14289 13141 14323 13175
rect 14323 13141 14332 13175
rect 14280 13132 14332 13141
rect 19892 13268 19944 13320
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 22100 13268 22152 13277
rect 24400 13311 24452 13320
rect 24400 13277 24409 13311
rect 24409 13277 24443 13311
rect 24443 13277 24452 13311
rect 24400 13268 24452 13277
rect 26240 13268 26292 13320
rect 17040 13243 17092 13252
rect 17040 13209 17049 13243
rect 17049 13209 17083 13243
rect 17083 13209 17092 13243
rect 17040 13200 17092 13209
rect 18604 13200 18656 13252
rect 25964 13200 26016 13252
rect 29460 13268 29512 13320
rect 30288 13311 30340 13320
rect 30288 13277 30297 13311
rect 30297 13277 30331 13311
rect 30331 13277 30340 13311
rect 30288 13268 30340 13277
rect 30840 13268 30892 13320
rect 32588 13336 32640 13388
rect 36912 13336 36964 13388
rect 36268 13268 36320 13320
rect 31024 13243 31076 13252
rect 31024 13209 31033 13243
rect 31033 13209 31067 13243
rect 31067 13209 31076 13243
rect 31024 13200 31076 13209
rect 31392 13200 31444 13252
rect 33692 13200 33744 13252
rect 35532 13200 35584 13252
rect 18788 13132 18840 13184
rect 25412 13132 25464 13184
rect 32220 13132 32272 13184
rect 33140 13132 33192 13184
rect 34796 13132 34848 13184
rect 40684 13336 40736 13388
rect 42616 13379 42668 13388
rect 42616 13345 42625 13379
rect 42625 13345 42659 13379
rect 42659 13345 42668 13379
rect 42616 13336 42668 13345
rect 40500 13311 40552 13320
rect 40500 13277 40509 13311
rect 40509 13277 40543 13311
rect 40543 13277 40552 13311
rect 40500 13268 40552 13277
rect 41144 13268 41196 13320
rect 41696 13268 41748 13320
rect 42800 13268 42852 13320
rect 43536 13311 43588 13320
rect 43536 13277 43545 13311
rect 43545 13277 43579 13311
rect 43579 13277 43588 13311
rect 43536 13268 43588 13277
rect 41328 13200 41380 13252
rect 42156 13243 42208 13252
rect 42156 13209 42165 13243
rect 42165 13209 42199 13243
rect 42199 13209 42208 13243
rect 43996 13472 44048 13524
rect 45468 13472 45520 13524
rect 52920 13472 52972 13524
rect 57980 13472 58032 13524
rect 45192 13336 45244 13388
rect 44824 13268 44876 13320
rect 42156 13200 42208 13209
rect 45376 13200 45428 13252
rect 45560 13311 45612 13320
rect 45560 13277 45569 13311
rect 45569 13277 45603 13311
rect 45603 13277 45612 13311
rect 46296 13311 46348 13320
rect 45560 13268 45612 13277
rect 46296 13277 46305 13311
rect 46305 13277 46339 13311
rect 46339 13277 46348 13311
rect 46296 13268 46348 13277
rect 47216 13311 47268 13320
rect 47216 13277 47225 13311
rect 47225 13277 47259 13311
rect 47259 13277 47268 13311
rect 47216 13268 47268 13277
rect 50620 13404 50672 13456
rect 51908 13379 51960 13388
rect 51908 13345 51917 13379
rect 51917 13345 51951 13379
rect 51951 13345 51960 13379
rect 51908 13336 51960 13345
rect 53380 13336 53432 13388
rect 56692 13379 56744 13388
rect 56692 13345 56701 13379
rect 56701 13345 56735 13379
rect 56735 13345 56744 13379
rect 56692 13336 56744 13345
rect 47492 13311 47544 13320
rect 47492 13277 47501 13311
rect 47501 13277 47535 13311
rect 47535 13277 47544 13311
rect 48228 13311 48280 13320
rect 47492 13268 47544 13277
rect 48228 13277 48237 13311
rect 48237 13277 48271 13311
rect 48271 13277 48280 13311
rect 48228 13268 48280 13277
rect 50344 13311 50396 13320
rect 50344 13277 50353 13311
rect 50353 13277 50387 13311
rect 50387 13277 50396 13311
rect 50344 13268 50396 13277
rect 50804 13311 50856 13320
rect 50804 13277 50813 13311
rect 50813 13277 50847 13311
rect 50847 13277 50856 13311
rect 50804 13268 50856 13277
rect 48780 13243 48832 13252
rect 38200 13132 38252 13184
rect 44916 13132 44968 13184
rect 47032 13175 47084 13184
rect 47032 13141 47041 13175
rect 47041 13141 47075 13175
rect 47075 13141 47084 13175
rect 47032 13132 47084 13141
rect 48780 13209 48789 13243
rect 48789 13209 48823 13243
rect 48823 13209 48832 13243
rect 48780 13200 48832 13209
rect 49792 13200 49844 13252
rect 51356 13268 51408 13320
rect 53564 13268 53616 13320
rect 55588 13268 55640 13320
rect 48320 13132 48372 13184
rect 49332 13132 49384 13184
rect 53196 13200 53248 13252
rect 57336 13200 57388 13252
rect 55312 13132 55364 13184
rect 15398 13030 15450 13082
rect 15462 13030 15514 13082
rect 15526 13030 15578 13082
rect 15590 13030 15642 13082
rect 15654 13030 15706 13082
rect 29846 13030 29898 13082
rect 29910 13030 29962 13082
rect 29974 13030 30026 13082
rect 30038 13030 30090 13082
rect 30102 13030 30154 13082
rect 44294 13030 44346 13082
rect 44358 13030 44410 13082
rect 44422 13030 44474 13082
rect 44486 13030 44538 13082
rect 44550 13030 44602 13082
rect 9680 12971 9732 12980
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 10048 12928 10100 12980
rect 16948 12928 17000 12980
rect 17960 12928 18012 12980
rect 18328 12928 18380 12980
rect 22468 12928 22520 12980
rect 23204 12928 23256 12980
rect 26516 12928 26568 12980
rect 30288 12928 30340 12980
rect 31116 12928 31168 12980
rect 10968 12903 11020 12912
rect 10968 12869 10977 12903
rect 10977 12869 11011 12903
rect 11011 12869 11020 12903
rect 10968 12860 11020 12869
rect 14372 12903 14424 12912
rect 14372 12869 14381 12903
rect 14381 12869 14415 12903
rect 14415 12869 14424 12903
rect 14372 12860 14424 12869
rect 17316 12903 17368 12912
rect 17316 12869 17325 12903
rect 17325 12869 17359 12903
rect 17359 12869 17368 12903
rect 17316 12860 17368 12869
rect 19984 12860 20036 12912
rect 23756 12860 23808 12912
rect 24216 12860 24268 12912
rect 7472 12792 7524 12844
rect 11152 12792 11204 12844
rect 11888 12792 11940 12844
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 12624 12835 12676 12844
rect 12624 12801 12633 12835
rect 12633 12801 12667 12835
rect 12667 12801 12676 12835
rect 12624 12792 12676 12801
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 19892 12835 19944 12844
rect 19892 12801 19901 12835
rect 19901 12801 19935 12835
rect 19935 12801 19944 12835
rect 19892 12792 19944 12801
rect 22100 12835 22152 12844
rect 7748 12767 7800 12776
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 13452 12724 13504 12776
rect 13728 12724 13780 12776
rect 17040 12724 17092 12776
rect 18604 12767 18656 12776
rect 15016 12656 15068 12708
rect 18604 12733 18613 12767
rect 18613 12733 18647 12767
rect 18647 12733 18656 12767
rect 18604 12724 18656 12733
rect 18972 12724 19024 12776
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 29460 12860 29512 12912
rect 29828 12903 29880 12912
rect 29828 12869 29837 12903
rect 29837 12869 29871 12903
rect 29871 12869 29880 12903
rect 29828 12860 29880 12869
rect 31208 12903 31260 12912
rect 31208 12869 31217 12903
rect 31217 12869 31251 12903
rect 31251 12869 31260 12903
rect 31208 12860 31260 12869
rect 35348 12928 35400 12980
rect 35532 12971 35584 12980
rect 35532 12937 35541 12971
rect 35541 12937 35575 12971
rect 35575 12937 35584 12971
rect 35532 12928 35584 12937
rect 39396 12928 39448 12980
rect 40960 12928 41012 12980
rect 41696 12928 41748 12980
rect 34796 12860 34848 12912
rect 48780 12928 48832 12980
rect 50436 12928 50488 12980
rect 33600 12792 33652 12844
rect 33784 12835 33836 12844
rect 33784 12801 33793 12835
rect 33793 12801 33827 12835
rect 33827 12801 33836 12835
rect 33784 12792 33836 12801
rect 35992 12835 36044 12844
rect 35992 12801 36001 12835
rect 36001 12801 36035 12835
rect 36035 12801 36044 12835
rect 35992 12792 36044 12801
rect 39396 12792 39448 12844
rect 40592 12792 40644 12844
rect 40960 12835 41012 12844
rect 40960 12801 40969 12835
rect 40969 12801 41003 12835
rect 41003 12801 41012 12835
rect 40960 12792 41012 12801
rect 43536 12792 43588 12844
rect 44732 12835 44784 12844
rect 44732 12801 44741 12835
rect 44741 12801 44775 12835
rect 44775 12801 44784 12835
rect 44732 12792 44784 12801
rect 44916 12835 44968 12844
rect 44916 12801 44925 12835
rect 44925 12801 44959 12835
rect 44959 12801 44968 12835
rect 44916 12792 44968 12801
rect 45192 12792 45244 12844
rect 23020 12724 23072 12776
rect 18144 12656 18196 12708
rect 7932 12631 7984 12640
rect 7932 12597 7941 12631
rect 7941 12597 7975 12631
rect 7975 12597 7984 12631
rect 7932 12588 7984 12597
rect 14280 12588 14332 12640
rect 17132 12588 17184 12640
rect 32220 12767 32272 12776
rect 23848 12631 23900 12640
rect 23848 12597 23857 12631
rect 23857 12597 23891 12631
rect 23891 12597 23900 12631
rect 23848 12588 23900 12597
rect 27620 12631 27672 12640
rect 27620 12597 27629 12631
rect 27629 12597 27663 12631
rect 27663 12597 27672 12631
rect 27620 12588 27672 12597
rect 32220 12733 32229 12767
rect 32229 12733 32263 12767
rect 32263 12733 32272 12767
rect 32220 12724 32272 12733
rect 33140 12767 33192 12776
rect 33140 12733 33149 12767
rect 33149 12733 33183 12767
rect 33183 12733 33192 12767
rect 33140 12724 33192 12733
rect 34060 12767 34112 12776
rect 34060 12733 34069 12767
rect 34069 12733 34103 12767
rect 34103 12733 34112 12767
rect 34060 12724 34112 12733
rect 35532 12724 35584 12776
rect 37464 12767 37516 12776
rect 37464 12733 37473 12767
rect 37473 12733 37507 12767
rect 37507 12733 37516 12767
rect 37464 12724 37516 12733
rect 40132 12767 40184 12776
rect 40132 12733 40141 12767
rect 40141 12733 40175 12767
rect 40175 12733 40184 12767
rect 40132 12724 40184 12733
rect 42156 12724 42208 12776
rect 45284 12724 45336 12776
rect 46756 12792 46808 12844
rect 48228 12792 48280 12844
rect 49332 12835 49384 12844
rect 49332 12801 49341 12835
rect 49341 12801 49375 12835
rect 49375 12801 49384 12835
rect 49332 12792 49384 12801
rect 50252 12860 50304 12912
rect 53196 12928 53248 12980
rect 53380 12971 53432 12980
rect 53380 12937 53389 12971
rect 53389 12937 53423 12971
rect 53423 12937 53432 12971
rect 53380 12928 53432 12937
rect 53564 12928 53616 12980
rect 51908 12860 51960 12912
rect 55680 12928 55732 12980
rect 58072 12971 58124 12980
rect 55312 12903 55364 12912
rect 55312 12869 55321 12903
rect 55321 12869 55355 12903
rect 55355 12869 55364 12903
rect 55312 12860 55364 12869
rect 50344 12792 50396 12844
rect 53012 12792 53064 12844
rect 55588 12835 55640 12844
rect 55588 12801 55597 12835
rect 55597 12801 55631 12835
rect 55631 12801 55640 12835
rect 55588 12792 55640 12801
rect 56048 12792 56100 12844
rect 57152 12835 57204 12844
rect 57152 12801 57161 12835
rect 57161 12801 57195 12835
rect 57195 12801 57204 12835
rect 57152 12792 57204 12801
rect 58072 12937 58081 12971
rect 58081 12937 58115 12971
rect 58115 12937 58124 12971
rect 58072 12928 58124 12937
rect 48136 12724 48188 12776
rect 49148 12767 49200 12776
rect 30932 12588 30984 12640
rect 31484 12588 31536 12640
rect 31668 12588 31720 12640
rect 33232 12656 33284 12708
rect 37648 12656 37700 12708
rect 41512 12656 41564 12708
rect 46940 12656 46992 12708
rect 48688 12699 48740 12708
rect 48688 12665 48697 12699
rect 48697 12665 48731 12699
rect 48731 12665 48740 12699
rect 48688 12656 48740 12665
rect 49148 12733 49157 12767
rect 49157 12733 49191 12767
rect 49191 12733 49200 12767
rect 49148 12724 49200 12733
rect 35440 12588 35492 12640
rect 38476 12588 38528 12640
rect 40132 12588 40184 12640
rect 45284 12588 45336 12640
rect 46480 12588 46532 12640
rect 48412 12588 48464 12640
rect 50804 12724 50856 12776
rect 53380 12767 53432 12776
rect 53380 12733 53389 12767
rect 53389 12733 53423 12767
rect 53423 12733 53432 12767
rect 53380 12724 53432 12733
rect 55680 12724 55732 12776
rect 53932 12656 53984 12708
rect 56600 12656 56652 12708
rect 52368 12588 52420 12640
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 8302 12486 8354 12538
rect 8366 12486 8418 12538
rect 8430 12486 8482 12538
rect 22622 12486 22674 12538
rect 22686 12486 22738 12538
rect 22750 12486 22802 12538
rect 22814 12486 22866 12538
rect 22878 12486 22930 12538
rect 37070 12486 37122 12538
rect 37134 12486 37186 12538
rect 37198 12486 37250 12538
rect 37262 12486 37314 12538
rect 37326 12486 37378 12538
rect 51518 12486 51570 12538
rect 51582 12486 51634 12538
rect 51646 12486 51698 12538
rect 51710 12486 51762 12538
rect 51774 12486 51826 12538
rect 10784 12384 10836 12436
rect 14740 12384 14792 12436
rect 16764 12384 16816 12436
rect 16856 12384 16908 12436
rect 19432 12384 19484 12436
rect 23756 12427 23808 12436
rect 23756 12393 23765 12427
rect 23765 12393 23799 12427
rect 23799 12393 23808 12427
rect 23756 12384 23808 12393
rect 13360 12248 13412 12300
rect 12624 12180 12676 12232
rect 13544 12180 13596 12232
rect 18236 12316 18288 12368
rect 18328 12316 18380 12368
rect 19524 12316 19576 12368
rect 20260 12316 20312 12368
rect 21364 12316 21416 12368
rect 30380 12384 30432 12436
rect 30656 12384 30708 12436
rect 31300 12384 31352 12436
rect 31392 12384 31444 12436
rect 33692 12384 33744 12436
rect 38752 12384 38804 12436
rect 41512 12384 41564 12436
rect 42156 12427 42208 12436
rect 42156 12393 42165 12427
rect 42165 12393 42199 12427
rect 42199 12393 42208 12427
rect 42156 12384 42208 12393
rect 29092 12316 29144 12368
rect 30288 12359 30340 12368
rect 30288 12325 30297 12359
rect 30297 12325 30331 12359
rect 30331 12325 30340 12359
rect 30288 12316 30340 12325
rect 31208 12316 31260 12368
rect 34060 12359 34112 12368
rect 18972 12180 19024 12232
rect 13084 12112 13136 12164
rect 16396 12155 16448 12164
rect 16396 12121 16405 12155
rect 16405 12121 16439 12155
rect 16439 12121 16448 12155
rect 16396 12112 16448 12121
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 16948 12044 17000 12096
rect 17132 12112 17184 12164
rect 21088 12180 21140 12232
rect 21824 12180 21876 12232
rect 24400 12248 24452 12300
rect 24584 12248 24636 12300
rect 28632 12248 28684 12300
rect 29552 12248 29604 12300
rect 33416 12248 33468 12300
rect 26148 12223 26200 12232
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 26424 12180 26476 12232
rect 26884 12223 26936 12232
rect 26884 12189 26893 12223
rect 26893 12189 26927 12223
rect 26927 12189 26936 12223
rect 26884 12180 26936 12189
rect 30656 12180 30708 12232
rect 31208 12223 31260 12232
rect 31208 12189 31217 12223
rect 31217 12189 31251 12223
rect 31251 12189 31260 12223
rect 31208 12180 31260 12189
rect 33692 12223 33744 12232
rect 22100 12112 22152 12164
rect 23204 12112 23256 12164
rect 25412 12112 25464 12164
rect 31024 12155 31076 12164
rect 31024 12121 31033 12155
rect 31033 12121 31067 12155
rect 31067 12121 31076 12155
rect 31024 12112 31076 12121
rect 33692 12189 33701 12223
rect 33701 12189 33735 12223
rect 33735 12189 33744 12223
rect 33692 12180 33744 12189
rect 34060 12325 34069 12359
rect 34069 12325 34103 12359
rect 34103 12325 34112 12359
rect 34060 12316 34112 12325
rect 36912 12316 36964 12368
rect 34796 12291 34848 12300
rect 34796 12257 34805 12291
rect 34805 12257 34839 12291
rect 34839 12257 34848 12291
rect 34796 12248 34848 12257
rect 35900 12248 35952 12300
rect 36360 12248 36412 12300
rect 34888 12223 34940 12232
rect 34520 12112 34572 12164
rect 34888 12189 34897 12223
rect 34897 12189 34931 12223
rect 34931 12189 34940 12223
rect 34888 12180 34940 12189
rect 36268 12180 36320 12232
rect 38108 12180 38160 12232
rect 39856 12316 39908 12368
rect 39764 12248 39816 12300
rect 40500 12248 40552 12300
rect 38476 12223 38528 12232
rect 38476 12189 38485 12223
rect 38485 12189 38519 12223
rect 38519 12189 38528 12223
rect 38476 12180 38528 12189
rect 38752 12223 38804 12232
rect 38752 12189 38761 12223
rect 38761 12189 38795 12223
rect 38795 12189 38804 12223
rect 39856 12223 39908 12232
rect 38752 12180 38804 12189
rect 39856 12189 39865 12223
rect 39865 12189 39899 12223
rect 39899 12189 39908 12223
rect 39856 12180 39908 12189
rect 40132 12223 40184 12232
rect 40132 12189 40141 12223
rect 40141 12189 40175 12223
rect 40175 12189 40184 12223
rect 40132 12180 40184 12189
rect 41144 12180 41196 12232
rect 41972 12223 42024 12232
rect 41972 12189 41981 12223
rect 41981 12189 42015 12223
rect 42015 12189 42024 12223
rect 41972 12180 42024 12189
rect 46296 12384 46348 12436
rect 48228 12384 48280 12436
rect 47032 12248 47084 12300
rect 48688 12291 48740 12300
rect 48688 12257 48697 12291
rect 48697 12257 48731 12291
rect 48731 12257 48740 12291
rect 48688 12248 48740 12257
rect 49976 12384 50028 12436
rect 50804 12384 50856 12436
rect 51908 12384 51960 12436
rect 53012 12384 53064 12436
rect 54116 12427 54168 12436
rect 54116 12393 54125 12427
rect 54125 12393 54159 12427
rect 54159 12393 54168 12427
rect 54116 12384 54168 12393
rect 54392 12427 54444 12436
rect 54392 12393 54401 12427
rect 54401 12393 54435 12427
rect 54435 12393 54444 12427
rect 54392 12384 54444 12393
rect 49700 12248 49752 12300
rect 53472 12248 53524 12300
rect 54300 12248 54352 12300
rect 54484 12248 54536 12300
rect 50436 12223 50488 12232
rect 39580 12112 39632 12164
rect 39764 12112 39816 12164
rect 42432 12112 42484 12164
rect 43628 12112 43680 12164
rect 18236 12044 18288 12096
rect 19432 12044 19484 12096
rect 20352 12087 20404 12096
rect 20352 12053 20361 12087
rect 20361 12053 20395 12087
rect 20395 12053 20404 12087
rect 20352 12044 20404 12053
rect 23756 12044 23808 12096
rect 24400 12044 24452 12096
rect 27620 12044 27672 12096
rect 28264 12044 28316 12096
rect 31576 12044 31628 12096
rect 33140 12044 33192 12096
rect 38292 12044 38344 12096
rect 40040 12044 40092 12096
rect 42156 12044 42208 12096
rect 44180 12044 44232 12096
rect 45376 12112 45428 12164
rect 48228 12112 48280 12164
rect 50436 12189 50445 12223
rect 50445 12189 50479 12223
rect 50479 12189 50488 12223
rect 50436 12180 50488 12189
rect 50804 12180 50856 12232
rect 52552 12112 52604 12164
rect 53380 12112 53432 12164
rect 53840 12112 53892 12164
rect 51080 12044 51132 12096
rect 53012 12044 53064 12096
rect 55680 12180 55732 12232
rect 56784 12155 56836 12164
rect 56784 12121 56793 12155
rect 56793 12121 56827 12155
rect 56827 12121 56836 12155
rect 56784 12112 56836 12121
rect 55312 12087 55364 12096
rect 55312 12053 55321 12087
rect 55321 12053 55355 12087
rect 55355 12053 55364 12087
rect 55312 12044 55364 12053
rect 15398 11942 15450 11994
rect 15462 11942 15514 11994
rect 15526 11942 15578 11994
rect 15590 11942 15642 11994
rect 15654 11942 15706 11994
rect 29846 11942 29898 11994
rect 29910 11942 29962 11994
rect 29974 11942 30026 11994
rect 30038 11942 30090 11994
rect 30102 11942 30154 11994
rect 44294 11942 44346 11994
rect 44358 11942 44410 11994
rect 44422 11942 44474 11994
rect 44486 11942 44538 11994
rect 44550 11942 44602 11994
rect 12256 11883 12308 11892
rect 12256 11849 12265 11883
rect 12265 11849 12299 11883
rect 12299 11849 12308 11883
rect 12256 11840 12308 11849
rect 13268 11883 13320 11892
rect 13268 11849 13277 11883
rect 13277 11849 13311 11883
rect 13311 11849 13320 11883
rect 13268 11840 13320 11849
rect 14832 11883 14884 11892
rect 14832 11849 14841 11883
rect 14841 11849 14875 11883
rect 14875 11849 14884 11883
rect 14832 11840 14884 11849
rect 17592 11840 17644 11892
rect 18696 11883 18748 11892
rect 18696 11849 18705 11883
rect 18705 11849 18739 11883
rect 18739 11849 18748 11883
rect 18696 11840 18748 11849
rect 19616 11883 19668 11892
rect 19616 11849 19625 11883
rect 19625 11849 19659 11883
rect 19659 11849 19668 11883
rect 19616 11840 19668 11849
rect 11980 11772 12032 11824
rect 16212 11772 16264 11824
rect 19524 11772 19576 11824
rect 23848 11840 23900 11892
rect 24768 11840 24820 11892
rect 26148 11840 26200 11892
rect 30656 11883 30708 11892
rect 30656 11849 30665 11883
rect 30665 11849 30699 11883
rect 30699 11849 30708 11883
rect 30656 11840 30708 11849
rect 30840 11840 30892 11892
rect 33416 11883 33468 11892
rect 33416 11849 33425 11883
rect 33425 11849 33459 11883
rect 33459 11849 33468 11883
rect 33416 11840 33468 11849
rect 34796 11840 34848 11892
rect 35532 11883 35584 11892
rect 35532 11849 35541 11883
rect 35541 11849 35575 11883
rect 35575 11849 35584 11883
rect 35532 11840 35584 11849
rect 38108 11840 38160 11892
rect 23756 11815 23808 11824
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 17040 11704 17092 11756
rect 17868 11704 17920 11756
rect 20260 11747 20312 11756
rect 20260 11713 20269 11747
rect 20269 11713 20303 11747
rect 20303 11713 20312 11747
rect 20260 11704 20312 11713
rect 16856 11636 16908 11688
rect 17408 11679 17460 11688
rect 17408 11645 17417 11679
rect 17417 11645 17451 11679
rect 17451 11645 17460 11679
rect 17408 11636 17460 11645
rect 19524 11636 19576 11688
rect 21364 11704 21416 11756
rect 21456 11704 21508 11756
rect 23756 11781 23765 11815
rect 23765 11781 23799 11815
rect 23799 11781 23808 11815
rect 23756 11772 23808 11781
rect 27068 11772 27120 11824
rect 28264 11815 28316 11824
rect 28264 11781 28273 11815
rect 28273 11781 28307 11815
rect 28307 11781 28316 11815
rect 28264 11772 28316 11781
rect 29552 11772 29604 11824
rect 30104 11772 30156 11824
rect 23480 11747 23532 11756
rect 23480 11713 23489 11747
rect 23489 11713 23523 11747
rect 23523 11713 23532 11747
rect 23480 11704 23532 11713
rect 30564 11747 30616 11756
rect 30564 11713 30573 11747
rect 30573 11713 30607 11747
rect 30607 11713 30616 11747
rect 30564 11704 30616 11713
rect 31208 11704 31260 11756
rect 31392 11747 31444 11756
rect 31392 11713 31401 11747
rect 31401 11713 31435 11747
rect 31435 11713 31444 11747
rect 31392 11704 31444 11713
rect 31576 11747 31628 11756
rect 31576 11713 31585 11747
rect 31585 11713 31619 11747
rect 31619 11713 31628 11747
rect 31576 11704 31628 11713
rect 31668 11704 31720 11756
rect 32496 11704 32548 11756
rect 33600 11747 33652 11756
rect 33600 11713 33609 11747
rect 33609 11713 33643 11747
rect 33643 11713 33652 11747
rect 33600 11704 33652 11713
rect 35992 11772 36044 11824
rect 37832 11772 37884 11824
rect 38568 11772 38620 11824
rect 34520 11747 34572 11756
rect 34520 11713 34529 11747
rect 34529 11713 34563 11747
rect 34563 11713 34572 11747
rect 34520 11704 34572 11713
rect 22468 11636 22520 11688
rect 24492 11636 24544 11688
rect 27804 11636 27856 11688
rect 29000 11636 29052 11688
rect 30196 11636 30248 11688
rect 31116 11636 31168 11688
rect 17684 11611 17736 11620
rect 17684 11577 17693 11611
rect 17693 11577 17727 11611
rect 17727 11577 17736 11611
rect 17684 11568 17736 11577
rect 15108 11500 15160 11552
rect 21088 11568 21140 11620
rect 30932 11611 30984 11620
rect 21364 11500 21416 11552
rect 30932 11577 30941 11611
rect 30941 11577 30975 11611
rect 30975 11577 30984 11611
rect 30932 11568 30984 11577
rect 32956 11636 33008 11688
rect 34888 11704 34940 11756
rect 35440 11747 35492 11756
rect 35440 11713 35449 11747
rect 35449 11713 35483 11747
rect 35483 11713 35492 11747
rect 35440 11704 35492 11713
rect 35900 11704 35952 11756
rect 32588 11500 32640 11552
rect 35348 11500 35400 11552
rect 36268 11543 36320 11552
rect 36268 11509 36277 11543
rect 36277 11509 36311 11543
rect 36311 11509 36320 11543
rect 36268 11500 36320 11509
rect 37648 11636 37700 11688
rect 38476 11636 38528 11688
rect 38844 11679 38896 11688
rect 38844 11645 38853 11679
rect 38853 11645 38887 11679
rect 38887 11645 38896 11679
rect 38844 11636 38896 11645
rect 39580 11679 39632 11688
rect 39580 11645 39589 11679
rect 39589 11645 39623 11679
rect 39623 11645 39632 11679
rect 39580 11636 39632 11645
rect 40684 11772 40736 11824
rect 41972 11840 42024 11892
rect 40592 11747 40644 11756
rect 40592 11713 40601 11747
rect 40601 11713 40635 11747
rect 40635 11713 40644 11747
rect 40592 11704 40644 11713
rect 40224 11568 40276 11620
rect 43812 11772 43864 11824
rect 44180 11772 44232 11824
rect 45376 11840 45428 11892
rect 45192 11772 45244 11824
rect 48320 11840 48372 11892
rect 49516 11840 49568 11892
rect 53932 11883 53984 11892
rect 53932 11849 53941 11883
rect 53941 11849 53975 11883
rect 53975 11849 53984 11883
rect 53932 11840 53984 11849
rect 56784 11840 56836 11892
rect 48228 11772 48280 11824
rect 40960 11704 41012 11756
rect 42432 11747 42484 11756
rect 42432 11713 42441 11747
rect 42441 11713 42475 11747
rect 42475 11713 42484 11747
rect 42432 11704 42484 11713
rect 43720 11704 43772 11756
rect 48136 11747 48188 11756
rect 48136 11713 48145 11747
rect 48145 11713 48179 11747
rect 48179 11713 48188 11747
rect 48136 11704 48188 11713
rect 43444 11636 43496 11688
rect 45100 11636 45152 11688
rect 38200 11500 38252 11552
rect 38292 11500 38344 11552
rect 42432 11500 42484 11552
rect 45376 11500 45428 11552
rect 45468 11500 45520 11552
rect 47860 11500 47912 11552
rect 49700 11704 49752 11756
rect 50896 11704 50948 11756
rect 48504 11636 48556 11688
rect 50436 11636 50488 11688
rect 51080 11679 51132 11688
rect 51080 11645 51089 11679
rect 51089 11645 51123 11679
rect 51123 11645 51132 11679
rect 51080 11636 51132 11645
rect 52000 11636 52052 11688
rect 53288 11704 53340 11756
rect 53932 11747 53984 11756
rect 53932 11713 53941 11747
rect 53941 11713 53975 11747
rect 53975 11713 53984 11747
rect 53932 11704 53984 11713
rect 54116 11704 54168 11756
rect 54944 11747 54996 11756
rect 54944 11713 54953 11747
rect 54953 11713 54987 11747
rect 54987 11713 54996 11747
rect 54944 11704 54996 11713
rect 55312 11704 55364 11756
rect 53012 11679 53064 11688
rect 53012 11645 53021 11679
rect 53021 11645 53055 11679
rect 53055 11645 53064 11679
rect 53012 11636 53064 11645
rect 53196 11636 53248 11688
rect 56140 11679 56192 11688
rect 56140 11645 56149 11679
rect 56149 11645 56183 11679
rect 56183 11645 56192 11679
rect 56140 11636 56192 11645
rect 52644 11568 52696 11620
rect 48964 11500 49016 11552
rect 50252 11543 50304 11552
rect 50252 11509 50261 11543
rect 50261 11509 50295 11543
rect 50295 11509 50304 11543
rect 50252 11500 50304 11509
rect 52092 11543 52144 11552
rect 52092 11509 52101 11543
rect 52101 11509 52135 11543
rect 52135 11509 52144 11543
rect 52092 11500 52144 11509
rect 53104 11500 53156 11552
rect 57796 11500 57848 11552
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 8302 11398 8354 11450
rect 8366 11398 8418 11450
rect 8430 11398 8482 11450
rect 22622 11398 22674 11450
rect 22686 11398 22738 11450
rect 22750 11398 22802 11450
rect 22814 11398 22866 11450
rect 22878 11398 22930 11450
rect 37070 11398 37122 11450
rect 37134 11398 37186 11450
rect 37198 11398 37250 11450
rect 37262 11398 37314 11450
rect 37326 11398 37378 11450
rect 51518 11398 51570 11450
rect 51582 11398 51634 11450
rect 51646 11398 51698 11450
rect 51710 11398 51762 11450
rect 51774 11398 51826 11450
rect 12808 11339 12860 11348
rect 12808 11305 12817 11339
rect 12817 11305 12851 11339
rect 12851 11305 12860 11339
rect 12808 11296 12860 11305
rect 13360 11296 13412 11348
rect 16672 11296 16724 11348
rect 18052 11296 18104 11348
rect 16028 11160 16080 11212
rect 19708 11160 19760 11212
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 20720 11160 20772 11212
rect 11888 11092 11940 11144
rect 15108 11135 15160 11144
rect 15108 11101 15117 11135
rect 15117 11101 15151 11135
rect 15151 11101 15160 11135
rect 15108 11092 15160 11101
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 17868 11092 17920 11144
rect 19524 11092 19576 11144
rect 16028 11067 16080 11076
rect 16028 11033 16037 11067
rect 16037 11033 16071 11067
rect 16071 11033 16080 11067
rect 16028 11024 16080 11033
rect 16580 11024 16632 11076
rect 21364 11228 21416 11280
rect 27344 11296 27396 11348
rect 28632 11339 28684 11348
rect 28632 11305 28641 11339
rect 28641 11305 28675 11339
rect 28675 11305 28684 11339
rect 28632 11296 28684 11305
rect 30932 11296 30984 11348
rect 31668 11296 31720 11348
rect 32956 11339 33008 11348
rect 32956 11305 32965 11339
rect 32965 11305 32999 11339
rect 32999 11305 33008 11339
rect 32956 11296 33008 11305
rect 34520 11296 34572 11348
rect 38844 11296 38896 11348
rect 42708 11296 42760 11348
rect 45100 11339 45152 11348
rect 45100 11305 45109 11339
rect 45109 11305 45143 11339
rect 45143 11305 45152 11339
rect 45100 11296 45152 11305
rect 45376 11296 45428 11348
rect 52092 11296 52144 11348
rect 53196 11339 53248 11348
rect 23848 11203 23900 11212
rect 23848 11169 23857 11203
rect 23857 11169 23891 11203
rect 23891 11169 23900 11203
rect 23848 11160 23900 11169
rect 24400 11092 24452 11144
rect 24676 11160 24728 11212
rect 24952 11092 25004 11144
rect 30564 11228 30616 11280
rect 30288 11160 30340 11212
rect 35348 11203 35400 11212
rect 35348 11169 35357 11203
rect 35357 11169 35391 11203
rect 35391 11169 35400 11203
rect 35348 11160 35400 11169
rect 35440 11160 35492 11212
rect 40132 11228 40184 11280
rect 40776 11228 40828 11280
rect 40960 11271 41012 11280
rect 40960 11237 40969 11271
rect 40969 11237 41003 11271
rect 41003 11237 41012 11271
rect 40960 11228 41012 11237
rect 43812 11228 43864 11280
rect 48504 11228 48556 11280
rect 36912 11160 36964 11212
rect 39948 11160 40000 11212
rect 22376 11067 22428 11076
rect 22376 11033 22385 11067
rect 22385 11033 22419 11067
rect 22419 11033 22428 11067
rect 22376 11024 22428 11033
rect 23848 11024 23900 11076
rect 25504 11024 25556 11076
rect 28172 11024 28224 11076
rect 30380 11092 30432 11144
rect 30104 11024 30156 11076
rect 31024 11092 31076 11144
rect 32588 11135 32640 11144
rect 32588 11101 32597 11135
rect 32597 11101 32631 11135
rect 32631 11101 32640 11135
rect 32588 11092 32640 11101
rect 35072 11135 35124 11144
rect 35072 11101 35081 11135
rect 35081 11101 35115 11135
rect 35115 11101 35124 11135
rect 35072 11092 35124 11101
rect 38108 11135 38160 11144
rect 38108 11101 38117 11135
rect 38117 11101 38151 11135
rect 38151 11101 38160 11135
rect 38108 11092 38160 11101
rect 38476 11092 38528 11144
rect 40040 11092 40092 11144
rect 33600 11024 33652 11076
rect 35440 11024 35492 11076
rect 36636 11024 36688 11076
rect 16212 10956 16264 11008
rect 17040 10956 17092 11008
rect 17408 10956 17460 11008
rect 17868 10956 17920 11008
rect 21916 10956 21968 11008
rect 26516 10956 26568 11008
rect 31668 10956 31720 11008
rect 32496 10956 32548 11008
rect 37280 11024 37332 11076
rect 38200 11024 38252 11076
rect 37924 10956 37976 11008
rect 41236 11160 41288 11212
rect 45284 11203 45336 11212
rect 45284 11169 45293 11203
rect 45293 11169 45327 11203
rect 45327 11169 45336 11203
rect 45284 11160 45336 11169
rect 44916 11092 44968 11144
rect 45468 11092 45520 11144
rect 48228 11160 48280 11212
rect 53196 11305 53205 11339
rect 53205 11305 53239 11339
rect 53239 11305 53248 11339
rect 53196 11296 53248 11305
rect 54944 11296 54996 11348
rect 57152 11296 57204 11348
rect 53288 11228 53340 11280
rect 56140 11160 56192 11212
rect 57796 11160 57848 11212
rect 47400 11135 47452 11144
rect 47400 11101 47409 11135
rect 47409 11101 47443 11135
rect 47443 11101 47452 11135
rect 47400 11092 47452 11101
rect 47860 11135 47912 11144
rect 47860 11101 47869 11135
rect 47869 11101 47903 11135
rect 47903 11101 47912 11135
rect 47860 11092 47912 11101
rect 48044 11092 48096 11144
rect 49700 11092 49752 11144
rect 49792 11092 49844 11144
rect 52644 11135 52696 11144
rect 52644 11101 52653 11135
rect 52653 11101 52687 11135
rect 52687 11101 52696 11135
rect 52644 11092 52696 11101
rect 53104 11135 53156 11144
rect 53104 11101 53113 11135
rect 53113 11101 53147 11135
rect 53147 11101 53156 11135
rect 53104 11092 53156 11101
rect 53932 11135 53984 11144
rect 42156 11024 42208 11076
rect 42432 11067 42484 11076
rect 42432 11033 42441 11067
rect 42441 11033 42475 11067
rect 42475 11033 42484 11067
rect 42432 11024 42484 11033
rect 50896 11024 50948 11076
rect 52000 11024 52052 11076
rect 53932 11101 53941 11135
rect 53941 11101 53975 11135
rect 53975 11101 53984 11135
rect 53932 11092 53984 11101
rect 56600 11024 56652 11076
rect 42340 10956 42392 11008
rect 43536 10999 43588 11008
rect 43536 10965 43545 10999
rect 43545 10965 43579 10999
rect 43579 10965 43588 10999
rect 43536 10956 43588 10965
rect 47400 10956 47452 11008
rect 48136 10956 48188 11008
rect 51908 10999 51960 11008
rect 51908 10965 51917 10999
rect 51917 10965 51951 10999
rect 51951 10965 51960 10999
rect 51908 10956 51960 10965
rect 15398 10854 15450 10906
rect 15462 10854 15514 10906
rect 15526 10854 15578 10906
rect 15590 10854 15642 10906
rect 15654 10854 15706 10906
rect 29846 10854 29898 10906
rect 29910 10854 29962 10906
rect 29974 10854 30026 10906
rect 30038 10854 30090 10906
rect 30102 10854 30154 10906
rect 44294 10854 44346 10906
rect 44358 10854 44410 10906
rect 44422 10854 44474 10906
rect 44486 10854 44538 10906
rect 44550 10854 44602 10906
rect 1860 10752 1912 10804
rect 16028 10752 16080 10804
rect 17960 10752 18012 10804
rect 18604 10752 18656 10804
rect 21180 10795 21232 10804
rect 16580 10684 16632 10736
rect 17592 10684 17644 10736
rect 1584 10616 1636 10668
rect 16212 10616 16264 10668
rect 17868 10684 17920 10736
rect 20444 10727 20496 10736
rect 20444 10693 20453 10727
rect 20453 10693 20487 10727
rect 20487 10693 20496 10727
rect 20444 10684 20496 10693
rect 19340 10616 19392 10668
rect 21180 10761 21189 10795
rect 21189 10761 21223 10795
rect 21223 10761 21232 10795
rect 21180 10752 21232 10761
rect 21916 10752 21968 10804
rect 22376 10684 22428 10736
rect 24492 10684 24544 10736
rect 21180 10616 21232 10668
rect 21916 10659 21968 10668
rect 21916 10625 21925 10659
rect 21925 10625 21959 10659
rect 21959 10625 21968 10659
rect 21916 10616 21968 10625
rect 25504 10616 25556 10668
rect 17684 10548 17736 10600
rect 20352 10548 20404 10600
rect 17040 10523 17092 10532
rect 17040 10489 17049 10523
rect 17049 10489 17083 10523
rect 17083 10489 17092 10523
rect 17040 10480 17092 10489
rect 23572 10548 23624 10600
rect 24492 10548 24544 10600
rect 29092 10684 29144 10736
rect 29184 10684 29236 10736
rect 31760 10616 31812 10668
rect 27160 10591 27212 10600
rect 27160 10557 27169 10591
rect 27169 10557 27203 10591
rect 27203 10557 27212 10591
rect 27160 10548 27212 10557
rect 29552 10591 29604 10600
rect 29552 10557 29561 10591
rect 29561 10557 29595 10591
rect 29595 10557 29604 10591
rect 29552 10548 29604 10557
rect 30196 10548 30248 10600
rect 30748 10591 30800 10600
rect 30748 10557 30757 10591
rect 30757 10557 30791 10591
rect 30791 10557 30800 10591
rect 30748 10548 30800 10557
rect 30380 10480 30432 10532
rect 30656 10480 30708 10532
rect 36636 10752 36688 10804
rect 38476 10752 38528 10804
rect 40960 10752 41012 10804
rect 42340 10752 42392 10804
rect 43444 10752 43496 10804
rect 52644 10752 52696 10804
rect 33784 10727 33836 10736
rect 33784 10693 33793 10727
rect 33793 10693 33827 10727
rect 33827 10693 33836 10727
rect 33784 10684 33836 10693
rect 38936 10684 38988 10736
rect 39212 10684 39264 10736
rect 37280 10616 37332 10668
rect 37740 10659 37792 10668
rect 37740 10625 37749 10659
rect 37749 10625 37783 10659
rect 37783 10625 37792 10659
rect 37740 10616 37792 10625
rect 37924 10616 37976 10668
rect 40316 10616 40368 10668
rect 42524 10616 42576 10668
rect 42616 10616 42668 10668
rect 48044 10684 48096 10736
rect 49700 10727 49752 10736
rect 43536 10616 43588 10668
rect 43812 10616 43864 10668
rect 49700 10693 49709 10727
rect 49709 10693 49743 10727
rect 49743 10693 49752 10727
rect 49700 10684 49752 10693
rect 51908 10684 51960 10736
rect 48964 10659 49016 10668
rect 48964 10625 48973 10659
rect 48973 10625 49007 10659
rect 49007 10625 49016 10659
rect 48964 10616 49016 10625
rect 37464 10480 37516 10532
rect 40040 10480 40092 10532
rect 41144 10480 41196 10532
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 20996 10412 21048 10464
rect 32588 10455 32640 10464
rect 32588 10421 32597 10455
rect 32597 10421 32631 10455
rect 32631 10421 32640 10455
rect 32588 10412 32640 10421
rect 39948 10412 40000 10464
rect 40224 10412 40276 10464
rect 43536 10412 43588 10464
rect 48136 10548 48188 10600
rect 49516 10659 49568 10668
rect 49516 10625 49525 10659
rect 49525 10625 49559 10659
rect 49559 10625 49568 10659
rect 49516 10616 49568 10625
rect 51356 10616 51408 10668
rect 52368 10616 52420 10668
rect 56048 10616 56100 10668
rect 51448 10523 51500 10532
rect 45376 10455 45428 10464
rect 45376 10421 45385 10455
rect 45385 10421 45419 10455
rect 45419 10421 45428 10455
rect 45376 10412 45428 10421
rect 45560 10412 45612 10464
rect 48044 10412 48096 10464
rect 51448 10489 51457 10523
rect 51457 10489 51491 10523
rect 51491 10489 51500 10523
rect 51448 10480 51500 10489
rect 54576 10480 54628 10532
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 8302 10310 8354 10362
rect 8366 10310 8418 10362
rect 8430 10310 8482 10362
rect 22622 10310 22674 10362
rect 22686 10310 22738 10362
rect 22750 10310 22802 10362
rect 22814 10310 22866 10362
rect 22878 10310 22930 10362
rect 37070 10310 37122 10362
rect 37134 10310 37186 10362
rect 37198 10310 37250 10362
rect 37262 10310 37314 10362
rect 37326 10310 37378 10362
rect 51518 10310 51570 10362
rect 51582 10310 51634 10362
rect 51646 10310 51698 10362
rect 51710 10310 51762 10362
rect 51774 10310 51826 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 16212 10251 16264 10260
rect 16212 10217 16221 10251
rect 16221 10217 16255 10251
rect 16255 10217 16264 10251
rect 16212 10208 16264 10217
rect 24584 10208 24636 10260
rect 16672 10140 16724 10192
rect 21180 10140 21232 10192
rect 30472 10208 30524 10260
rect 30656 10251 30708 10260
rect 30656 10217 30665 10251
rect 30665 10217 30699 10251
rect 30699 10217 30708 10251
rect 30656 10208 30708 10217
rect 31024 10208 31076 10260
rect 31484 10251 31536 10260
rect 31484 10217 31493 10251
rect 31493 10217 31527 10251
rect 31527 10217 31536 10251
rect 31484 10208 31536 10217
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 18144 10072 18196 10081
rect 20260 10004 20312 10056
rect 19340 9936 19392 9988
rect 26240 10072 26292 10124
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 27712 10140 27764 10192
rect 28264 10140 28316 10192
rect 27160 10115 27212 10124
rect 27160 10081 27169 10115
rect 27169 10081 27203 10115
rect 27203 10081 27212 10115
rect 27160 10072 27212 10081
rect 28724 10072 28776 10124
rect 29368 10140 29420 10192
rect 30840 10072 30892 10124
rect 31668 10140 31720 10192
rect 32588 10208 32640 10260
rect 40592 10251 40644 10260
rect 40592 10217 40601 10251
rect 40601 10217 40635 10251
rect 40635 10217 40644 10251
rect 40592 10208 40644 10217
rect 40776 10208 40828 10260
rect 45560 10251 45612 10260
rect 45560 10217 45569 10251
rect 45569 10217 45603 10251
rect 45603 10217 45612 10251
rect 45560 10208 45612 10217
rect 48044 10208 48096 10260
rect 33324 10140 33376 10192
rect 41420 10140 41472 10192
rect 31852 10072 31904 10124
rect 21088 10004 21140 10056
rect 22100 10047 22152 10056
rect 22100 10013 22109 10047
rect 22109 10013 22143 10047
rect 22143 10013 22152 10047
rect 22100 10004 22152 10013
rect 13820 9868 13872 9920
rect 15752 9868 15804 9920
rect 18604 9868 18656 9920
rect 18788 9868 18840 9920
rect 20260 9911 20312 9920
rect 20260 9877 20269 9911
rect 20269 9877 20303 9911
rect 20303 9877 20312 9911
rect 20260 9868 20312 9877
rect 24676 9936 24728 9988
rect 30472 10047 30524 10056
rect 30472 10013 30481 10047
rect 30481 10013 30515 10047
rect 30515 10013 30524 10047
rect 30472 10004 30524 10013
rect 31760 10004 31812 10056
rect 33692 10072 33744 10124
rect 34704 10115 34756 10124
rect 34704 10081 34713 10115
rect 34713 10081 34747 10115
rect 34747 10081 34756 10115
rect 34704 10072 34756 10081
rect 35072 10072 35124 10124
rect 36912 10115 36964 10124
rect 36912 10081 36921 10115
rect 36921 10081 36955 10115
rect 36955 10081 36964 10115
rect 36912 10072 36964 10081
rect 38660 10115 38712 10124
rect 38660 10081 38669 10115
rect 38669 10081 38703 10115
rect 38703 10081 38712 10115
rect 38660 10072 38712 10081
rect 40040 10115 40092 10124
rect 40040 10081 40049 10115
rect 40049 10081 40083 10115
rect 40083 10081 40092 10115
rect 40040 10072 40092 10081
rect 40224 10072 40276 10124
rect 41236 10072 41288 10124
rect 51080 10115 51132 10124
rect 51080 10081 51089 10115
rect 51089 10081 51123 10115
rect 51123 10081 51132 10115
rect 53932 10208 53984 10260
rect 55404 10140 55456 10192
rect 51080 10072 51132 10081
rect 39120 10047 39172 10056
rect 28724 9936 28776 9988
rect 31668 9979 31720 9988
rect 31668 9945 31677 9979
rect 31677 9945 31711 9979
rect 31711 9945 31720 9979
rect 31668 9936 31720 9945
rect 26424 9868 26476 9920
rect 30840 9868 30892 9920
rect 33140 9936 33192 9988
rect 34612 9936 34664 9988
rect 34336 9868 34388 9920
rect 39120 10013 39129 10047
rect 39129 10013 39163 10047
rect 39163 10013 39172 10047
rect 39120 10004 39172 10013
rect 39304 10047 39356 10056
rect 39304 10013 39313 10047
rect 39313 10013 39347 10047
rect 39347 10013 39356 10047
rect 39304 10004 39356 10013
rect 51356 10047 51408 10056
rect 51356 10013 51365 10047
rect 51365 10013 51399 10047
rect 51399 10013 51408 10047
rect 51356 10004 51408 10013
rect 52368 10047 52420 10056
rect 52368 10013 52377 10047
rect 52377 10013 52411 10047
rect 52411 10013 52420 10047
rect 52368 10004 52420 10013
rect 36268 9936 36320 9988
rect 38200 9936 38252 9988
rect 38476 9936 38528 9988
rect 42524 9936 42576 9988
rect 42708 9936 42760 9988
rect 45468 9979 45520 9988
rect 45468 9945 45477 9979
rect 45477 9945 45511 9979
rect 45511 9945 45520 9979
rect 45468 9936 45520 9945
rect 51908 9936 51960 9988
rect 55128 10072 55180 10124
rect 56600 10072 56652 10124
rect 57336 10072 57388 10124
rect 52644 10047 52696 10056
rect 52644 10013 52653 10047
rect 52653 10013 52687 10047
rect 52687 10013 52696 10047
rect 52644 10004 52696 10013
rect 57520 9936 57572 9988
rect 38108 9868 38160 9920
rect 40132 9911 40184 9920
rect 40132 9877 40141 9911
rect 40141 9877 40175 9911
rect 40175 9877 40184 9911
rect 40132 9868 40184 9877
rect 41144 9868 41196 9920
rect 41236 9868 41288 9920
rect 44180 9868 44232 9920
rect 15398 9766 15450 9818
rect 15462 9766 15514 9818
rect 15526 9766 15578 9818
rect 15590 9766 15642 9818
rect 15654 9766 15706 9818
rect 29846 9766 29898 9818
rect 29910 9766 29962 9818
rect 29974 9766 30026 9818
rect 30038 9766 30090 9818
rect 30102 9766 30154 9818
rect 44294 9766 44346 9818
rect 44358 9766 44410 9818
rect 44422 9766 44474 9818
rect 44486 9766 44538 9818
rect 44550 9766 44602 9818
rect 17592 9664 17644 9716
rect 20260 9664 20312 9716
rect 20444 9664 20496 9716
rect 21916 9664 21968 9716
rect 20720 9639 20772 9648
rect 20720 9605 20729 9639
rect 20729 9605 20763 9639
rect 20763 9605 20772 9639
rect 20720 9596 20772 9605
rect 22468 9596 22520 9648
rect 23848 9528 23900 9580
rect 18420 9503 18472 9512
rect 3240 9324 3292 9376
rect 17776 9392 17828 9444
rect 16304 9324 16356 9376
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 18696 9503 18748 9512
rect 18696 9469 18705 9503
rect 18705 9469 18739 9503
rect 18739 9469 18748 9503
rect 18696 9460 18748 9469
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 30656 9664 30708 9716
rect 34612 9664 34664 9716
rect 28448 9596 28500 9648
rect 29276 9596 29328 9648
rect 36268 9664 36320 9716
rect 40132 9664 40184 9716
rect 42616 9664 42668 9716
rect 43536 9707 43588 9716
rect 43536 9673 43545 9707
rect 43545 9673 43579 9707
rect 43579 9673 43588 9707
rect 43536 9664 43588 9673
rect 38384 9639 38436 9648
rect 38384 9605 38393 9639
rect 38393 9605 38427 9639
rect 38427 9605 38436 9639
rect 38384 9596 38436 9605
rect 40040 9596 40092 9648
rect 41236 9596 41288 9648
rect 44824 9596 44876 9648
rect 49792 9664 49844 9716
rect 57520 9664 57572 9716
rect 31944 9528 31996 9580
rect 33692 9571 33744 9580
rect 33692 9537 33701 9571
rect 33701 9537 33735 9571
rect 33735 9537 33744 9571
rect 33692 9528 33744 9537
rect 35992 9528 36044 9580
rect 36912 9528 36964 9580
rect 41328 9528 41380 9580
rect 44732 9528 44784 9580
rect 45468 9528 45520 9580
rect 48228 9528 48280 9580
rect 51448 9596 51500 9648
rect 52644 9596 52696 9648
rect 54576 9639 54628 9648
rect 54576 9605 54585 9639
rect 54585 9605 54619 9639
rect 54619 9605 54628 9639
rect 54576 9596 54628 9605
rect 56600 9596 56652 9648
rect 50252 9528 50304 9580
rect 54300 9571 54352 9580
rect 54300 9537 54309 9571
rect 54309 9537 54343 9571
rect 54343 9537 54352 9571
rect 54300 9528 54352 9537
rect 28080 9460 28132 9512
rect 30564 9460 30616 9512
rect 30656 9503 30708 9512
rect 30656 9469 30665 9503
rect 30665 9469 30699 9503
rect 30699 9469 30708 9503
rect 33968 9503 34020 9512
rect 30656 9460 30708 9469
rect 33968 9469 33977 9503
rect 33977 9469 34011 9503
rect 34011 9469 34020 9503
rect 33968 9460 34020 9469
rect 38844 9460 38896 9512
rect 40960 9460 41012 9512
rect 48320 9460 48372 9512
rect 27988 9392 28040 9444
rect 31760 9392 31812 9444
rect 20260 9324 20312 9376
rect 27252 9324 27304 9376
rect 28172 9324 28224 9376
rect 30196 9324 30248 9376
rect 30380 9324 30432 9376
rect 33692 9392 33744 9444
rect 35072 9392 35124 9444
rect 35900 9392 35952 9444
rect 39304 9392 39356 9444
rect 33324 9324 33376 9376
rect 38936 9324 38988 9376
rect 39764 9324 39816 9376
rect 46940 9392 46992 9444
rect 51080 9460 51132 9512
rect 56048 9503 56100 9512
rect 56048 9469 56057 9503
rect 56057 9469 56091 9503
rect 56091 9469 56100 9503
rect 56048 9460 56100 9469
rect 40868 9324 40920 9376
rect 41052 9324 41104 9376
rect 42892 9367 42944 9376
rect 42892 9333 42901 9367
rect 42901 9333 42935 9367
rect 42935 9333 42944 9367
rect 42892 9324 42944 9333
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 8302 9222 8354 9274
rect 8366 9222 8418 9274
rect 8430 9222 8482 9274
rect 22622 9222 22674 9274
rect 22686 9222 22738 9274
rect 22750 9222 22802 9274
rect 22814 9222 22866 9274
rect 22878 9222 22930 9274
rect 37070 9222 37122 9274
rect 37134 9222 37186 9274
rect 37198 9222 37250 9274
rect 37262 9222 37314 9274
rect 37326 9222 37378 9274
rect 51518 9222 51570 9274
rect 51582 9222 51634 9274
rect 51646 9222 51698 9274
rect 51710 9222 51762 9274
rect 51774 9222 51826 9274
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 18696 9120 18748 9172
rect 19892 9120 19944 9172
rect 20996 9163 21048 9172
rect 20996 9129 21005 9163
rect 21005 9129 21039 9163
rect 21039 9129 21048 9163
rect 20996 9120 21048 9129
rect 33968 9120 34020 9172
rect 34152 9120 34204 9172
rect 20260 9095 20312 9104
rect 20260 9061 20269 9095
rect 20269 9061 20303 9095
rect 20303 9061 20312 9095
rect 20260 9052 20312 9061
rect 27252 9052 27304 9104
rect 26424 8959 26476 8968
rect 26424 8925 26433 8959
rect 26433 8925 26467 8959
rect 26467 8925 26476 8959
rect 26424 8916 26476 8925
rect 27252 8959 27304 8968
rect 27252 8925 27261 8959
rect 27261 8925 27295 8959
rect 27295 8925 27304 8959
rect 27252 8916 27304 8925
rect 29368 8984 29420 9036
rect 29644 9027 29696 9036
rect 29644 8993 29653 9027
rect 29653 8993 29687 9027
rect 29687 8993 29696 9027
rect 29644 8984 29696 8993
rect 17132 8891 17184 8900
rect 17132 8857 17141 8891
rect 17141 8857 17175 8891
rect 17175 8857 17184 8891
rect 17132 8848 17184 8857
rect 17592 8848 17644 8900
rect 19984 8891 20036 8900
rect 19984 8857 19993 8891
rect 19993 8857 20027 8891
rect 20027 8857 20036 8891
rect 19984 8848 20036 8857
rect 1676 8780 1728 8832
rect 16304 8823 16356 8832
rect 16304 8789 16313 8823
rect 16313 8789 16347 8823
rect 16347 8789 16356 8823
rect 16304 8780 16356 8789
rect 20444 8823 20496 8832
rect 20444 8789 20453 8823
rect 20453 8789 20487 8823
rect 20487 8789 20496 8823
rect 20444 8780 20496 8789
rect 21180 8780 21232 8832
rect 28172 8959 28224 8968
rect 28172 8925 28181 8959
rect 28181 8925 28215 8959
rect 28215 8925 28224 8959
rect 29736 8959 29788 8968
rect 28172 8916 28224 8925
rect 29736 8925 29745 8959
rect 29745 8925 29779 8959
rect 29779 8925 29788 8959
rect 29736 8916 29788 8925
rect 30472 8984 30524 9036
rect 31576 9027 31628 9036
rect 31576 8993 31585 9027
rect 31585 8993 31619 9027
rect 31619 8993 31628 9027
rect 31576 8984 31628 8993
rect 33692 9052 33744 9104
rect 35072 9052 35124 9104
rect 34888 8984 34940 9036
rect 31944 8916 31996 8968
rect 32404 8959 32456 8968
rect 32404 8925 32413 8959
rect 32413 8925 32447 8959
rect 32447 8925 32456 8959
rect 32404 8916 32456 8925
rect 38568 9120 38620 9172
rect 40868 9120 40920 9172
rect 38660 9052 38712 9104
rect 38752 9052 38804 9104
rect 28724 8848 28776 8900
rect 31484 8848 31536 8900
rect 32680 8891 32732 8900
rect 32680 8857 32689 8891
rect 32689 8857 32723 8891
rect 32723 8857 32732 8891
rect 32680 8848 32732 8857
rect 34336 8848 34388 8900
rect 34428 8848 34480 8900
rect 35440 8891 35492 8900
rect 35440 8857 35449 8891
rect 35449 8857 35483 8891
rect 35483 8857 35492 8891
rect 35440 8848 35492 8857
rect 38200 8984 38252 9036
rect 39120 8984 39172 9036
rect 41328 9120 41380 9172
rect 42892 9120 42944 9172
rect 48228 9163 48280 9172
rect 48228 9129 48237 9163
rect 48237 9129 48271 9163
rect 48271 9129 48280 9163
rect 48228 9120 48280 9129
rect 50988 9120 51040 9172
rect 55128 9120 55180 9172
rect 45560 9052 45612 9104
rect 42340 8984 42392 9036
rect 46204 8984 46256 9036
rect 57336 9027 57388 9036
rect 57336 8993 57345 9027
rect 57345 8993 57379 9027
rect 57379 8993 57388 9027
rect 57336 8984 57388 8993
rect 38016 8916 38068 8968
rect 38292 8916 38344 8968
rect 38660 8916 38712 8968
rect 38844 8959 38896 8968
rect 38844 8925 38853 8959
rect 38853 8925 38887 8959
rect 38887 8925 38896 8959
rect 39028 8959 39080 8968
rect 38844 8916 38896 8925
rect 39028 8925 39037 8959
rect 39037 8925 39071 8959
rect 39071 8925 39080 8959
rect 39028 8916 39080 8925
rect 40040 8959 40092 8968
rect 40040 8925 40049 8959
rect 40049 8925 40083 8959
rect 40083 8925 40092 8959
rect 40040 8916 40092 8925
rect 40316 8959 40368 8968
rect 40316 8925 40325 8959
rect 40325 8925 40359 8959
rect 40359 8925 40368 8959
rect 40316 8916 40368 8925
rect 44088 8916 44140 8968
rect 45100 8916 45152 8968
rect 39304 8848 39356 8900
rect 42432 8848 42484 8900
rect 44180 8848 44232 8900
rect 31392 8780 31444 8832
rect 32312 8780 32364 8832
rect 34244 8780 34296 8832
rect 35072 8780 35124 8832
rect 36912 8780 36964 8832
rect 37740 8780 37792 8832
rect 39120 8780 39172 8832
rect 42892 8780 42944 8832
rect 45928 8848 45980 8900
rect 45192 8823 45244 8832
rect 45192 8789 45201 8823
rect 45201 8789 45235 8823
rect 45235 8789 45244 8823
rect 45192 8780 45244 8789
rect 45376 8780 45428 8832
rect 46388 8780 46440 8832
rect 47676 8780 47728 8832
rect 55588 8823 55640 8832
rect 55588 8789 55597 8823
rect 55597 8789 55631 8823
rect 55631 8789 55640 8823
rect 55588 8780 55640 8789
rect 56600 8848 56652 8900
rect 57796 8780 57848 8832
rect 15398 8678 15450 8730
rect 15462 8678 15514 8730
rect 15526 8678 15578 8730
rect 15590 8678 15642 8730
rect 15654 8678 15706 8730
rect 29846 8678 29898 8730
rect 29910 8678 29962 8730
rect 29974 8678 30026 8730
rect 30038 8678 30090 8730
rect 30102 8678 30154 8730
rect 44294 8678 44346 8730
rect 44358 8678 44410 8730
rect 44422 8678 44474 8730
rect 44486 8678 44538 8730
rect 44550 8678 44602 8730
rect 17132 8576 17184 8628
rect 19984 8576 20036 8628
rect 26424 8576 26476 8628
rect 28724 8576 28776 8628
rect 29368 8619 29420 8628
rect 20260 8508 20312 8560
rect 18788 8440 18840 8492
rect 28172 8508 28224 8560
rect 29368 8585 29377 8619
rect 29377 8585 29411 8619
rect 29411 8585 29420 8619
rect 29368 8576 29420 8585
rect 29644 8576 29696 8628
rect 31484 8619 31536 8628
rect 31484 8585 31493 8619
rect 31493 8585 31527 8619
rect 31527 8585 31536 8619
rect 31484 8576 31536 8585
rect 32680 8619 32732 8628
rect 32680 8585 32689 8619
rect 32689 8585 32723 8619
rect 32723 8585 32732 8619
rect 32680 8576 32732 8585
rect 32772 8576 32824 8628
rect 33048 8576 33100 8628
rect 34336 8576 34388 8628
rect 28448 8483 28500 8492
rect 28448 8449 28457 8483
rect 28457 8449 28491 8483
rect 28491 8449 28500 8483
rect 28448 8440 28500 8449
rect 30288 8440 30340 8492
rect 32128 8508 32180 8560
rect 35992 8576 36044 8628
rect 38476 8576 38528 8628
rect 39948 8576 40000 8628
rect 40960 8619 41012 8628
rect 35440 8508 35492 8560
rect 30840 8483 30892 8492
rect 19984 8304 20036 8356
rect 20536 8304 20588 8356
rect 29644 8304 29696 8356
rect 21180 8236 21232 8288
rect 27712 8236 27764 8288
rect 28816 8236 28868 8288
rect 30472 8304 30524 8356
rect 30840 8449 30849 8483
rect 30849 8449 30883 8483
rect 30883 8449 30892 8483
rect 30840 8440 30892 8449
rect 30932 8483 30984 8492
rect 30932 8449 30941 8483
rect 30941 8449 30975 8483
rect 30975 8449 30984 8483
rect 32312 8483 32364 8492
rect 30932 8440 30984 8449
rect 30748 8372 30800 8424
rect 32312 8449 32321 8483
rect 32321 8449 32355 8483
rect 32355 8449 32364 8483
rect 32312 8440 32364 8449
rect 39120 8508 39172 8560
rect 39304 8508 39356 8560
rect 32036 8372 32088 8424
rect 32220 8415 32272 8424
rect 32220 8381 32229 8415
rect 32229 8381 32263 8415
rect 32263 8381 32272 8415
rect 32220 8372 32272 8381
rect 32404 8372 32456 8424
rect 34888 8415 34940 8424
rect 34888 8381 34897 8415
rect 34897 8381 34931 8415
rect 34931 8381 34940 8415
rect 34888 8372 34940 8381
rect 31760 8304 31812 8356
rect 36912 8440 36964 8492
rect 38568 8483 38620 8492
rect 38384 8415 38436 8424
rect 38384 8381 38393 8415
rect 38393 8381 38427 8415
rect 38427 8381 38436 8415
rect 38384 8372 38436 8381
rect 38568 8449 38597 8483
rect 38597 8449 38620 8483
rect 38568 8440 38620 8449
rect 39856 8483 39908 8492
rect 39856 8449 39865 8483
rect 39865 8449 39899 8483
rect 39899 8449 39908 8483
rect 39856 8440 39908 8449
rect 40960 8585 40969 8619
rect 40969 8585 41003 8619
rect 41003 8585 41012 8619
rect 40960 8576 41012 8585
rect 42892 8576 42944 8628
rect 44732 8576 44784 8628
rect 45100 8576 45152 8628
rect 45560 8576 45612 8628
rect 46204 8619 46256 8628
rect 46204 8585 46213 8619
rect 46213 8585 46247 8619
rect 46247 8585 46256 8619
rect 46204 8576 46256 8585
rect 55404 8619 55456 8628
rect 55404 8585 55413 8619
rect 55413 8585 55447 8619
rect 55447 8585 55456 8619
rect 55404 8576 55456 8585
rect 39672 8372 39724 8424
rect 39948 8415 40000 8424
rect 39948 8381 39957 8415
rect 39957 8381 39991 8415
rect 39991 8381 40000 8415
rect 41604 8483 41656 8492
rect 41604 8449 41613 8483
rect 41613 8449 41647 8483
rect 41647 8449 41656 8483
rect 41604 8440 41656 8449
rect 44364 8483 44416 8492
rect 44364 8449 44373 8483
rect 44373 8449 44407 8483
rect 44407 8449 44416 8483
rect 44364 8440 44416 8449
rect 44640 8483 44692 8492
rect 44640 8449 44649 8483
rect 44649 8449 44683 8483
rect 44683 8449 44692 8483
rect 44640 8440 44692 8449
rect 45100 8440 45152 8492
rect 45376 8483 45428 8492
rect 45376 8449 45385 8483
rect 45385 8449 45419 8483
rect 45419 8449 45428 8483
rect 45376 8440 45428 8449
rect 46388 8483 46440 8492
rect 46388 8449 46397 8483
rect 46397 8449 46431 8483
rect 46431 8449 46440 8483
rect 46388 8440 46440 8449
rect 46572 8483 46624 8492
rect 46572 8449 46581 8483
rect 46581 8449 46615 8483
rect 46615 8449 46624 8483
rect 46572 8440 46624 8449
rect 47308 8440 47360 8492
rect 39948 8372 40000 8381
rect 40960 8415 41012 8424
rect 40960 8381 40969 8415
rect 40969 8381 41003 8415
rect 41003 8381 41012 8415
rect 40960 8372 41012 8381
rect 42616 8372 42668 8424
rect 31576 8236 31628 8288
rect 34152 8236 34204 8288
rect 34520 8236 34572 8288
rect 38476 8304 38528 8356
rect 39764 8304 39816 8356
rect 41420 8347 41472 8356
rect 41420 8313 41429 8347
rect 41429 8313 41463 8347
rect 41463 8313 41472 8347
rect 41420 8304 41472 8313
rect 37464 8236 37516 8288
rect 39948 8236 40000 8288
rect 40408 8236 40460 8288
rect 40500 8236 40552 8288
rect 41328 8236 41380 8288
rect 43076 8279 43128 8288
rect 43076 8245 43085 8279
rect 43085 8245 43119 8279
rect 43119 8245 43128 8279
rect 43076 8236 43128 8245
rect 44272 8236 44324 8288
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 8302 8134 8354 8186
rect 8366 8134 8418 8186
rect 8430 8134 8482 8186
rect 22622 8134 22674 8186
rect 22686 8134 22738 8186
rect 22750 8134 22802 8186
rect 22814 8134 22866 8186
rect 22878 8134 22930 8186
rect 37070 8134 37122 8186
rect 37134 8134 37186 8186
rect 37198 8134 37250 8186
rect 37262 8134 37314 8186
rect 37326 8134 37378 8186
rect 51518 8134 51570 8186
rect 51582 8134 51634 8186
rect 51646 8134 51698 8186
rect 51710 8134 51762 8186
rect 51774 8134 51826 8186
rect 21180 8075 21232 8084
rect 21180 8041 21189 8075
rect 21189 8041 21223 8075
rect 21223 8041 21232 8075
rect 21180 8032 21232 8041
rect 26424 8032 26476 8084
rect 28172 8032 28224 8084
rect 30840 8075 30892 8084
rect 30840 8041 30849 8075
rect 30849 8041 30883 8075
rect 30883 8041 30892 8075
rect 30840 8032 30892 8041
rect 32220 8032 32272 8084
rect 33048 8032 33100 8084
rect 30932 7964 30984 8016
rect 31668 8007 31720 8016
rect 31668 7973 31677 8007
rect 31677 7973 31711 8007
rect 31711 7973 31720 8007
rect 31668 7964 31720 7973
rect 31760 7964 31812 8016
rect 36912 8032 36964 8084
rect 27804 7896 27856 7948
rect 28632 7896 28684 7948
rect 29460 7896 29512 7948
rect 30564 7939 30616 7948
rect 30564 7905 30573 7939
rect 30573 7905 30607 7939
rect 30607 7905 30616 7939
rect 30564 7896 30616 7905
rect 20444 7828 20496 7880
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 28080 7871 28132 7880
rect 20536 7828 20588 7837
rect 28080 7837 28089 7871
rect 28089 7837 28123 7871
rect 28123 7837 28132 7871
rect 28080 7828 28132 7837
rect 28724 7871 28776 7880
rect 28724 7837 28733 7871
rect 28733 7837 28767 7871
rect 28767 7837 28776 7871
rect 28724 7828 28776 7837
rect 29736 7828 29788 7880
rect 32220 7896 32272 7948
rect 33048 7896 33100 7948
rect 34244 7896 34296 7948
rect 34704 7939 34756 7948
rect 34704 7905 34713 7939
rect 34713 7905 34747 7939
rect 34747 7905 34756 7939
rect 34704 7896 34756 7905
rect 37464 7964 37516 8016
rect 38476 7939 38528 7948
rect 38476 7905 38485 7939
rect 38485 7905 38519 7939
rect 38519 7905 38528 7939
rect 38476 7896 38528 7905
rect 40224 8032 40276 8084
rect 44364 8032 44416 8084
rect 47308 8075 47360 8084
rect 47308 8041 47317 8075
rect 47317 8041 47351 8075
rect 47351 8041 47360 8075
rect 47308 8032 47360 8041
rect 39856 7964 39908 8016
rect 40040 7896 40092 7948
rect 42340 7939 42392 7948
rect 42340 7905 42349 7939
rect 42349 7905 42383 7939
rect 42383 7905 42392 7939
rect 42340 7896 42392 7905
rect 57796 7964 57848 8016
rect 32036 7828 32088 7880
rect 32496 7828 32548 7880
rect 33692 7871 33744 7880
rect 33692 7837 33701 7871
rect 33701 7837 33735 7871
rect 33735 7837 33744 7871
rect 33692 7828 33744 7837
rect 34520 7828 34572 7880
rect 45376 7871 45428 7880
rect 45376 7837 45385 7871
rect 45385 7837 45419 7871
rect 45419 7837 45428 7871
rect 45376 7828 45428 7837
rect 46388 7896 46440 7948
rect 46296 7828 46348 7880
rect 27804 7803 27856 7812
rect 27804 7769 27813 7803
rect 27813 7769 27847 7803
rect 27847 7769 27856 7803
rect 27804 7760 27856 7769
rect 31300 7760 31352 7812
rect 20904 7692 20956 7744
rect 28448 7692 28500 7744
rect 29092 7692 29144 7744
rect 31576 7760 31628 7812
rect 32128 7760 32180 7812
rect 32680 7760 32732 7812
rect 35992 7760 36044 7812
rect 38016 7760 38068 7812
rect 38476 7760 38528 7812
rect 40408 7803 40460 7812
rect 40408 7769 40417 7803
rect 40417 7769 40451 7803
rect 40451 7769 40460 7803
rect 40408 7760 40460 7769
rect 41696 7760 41748 7812
rect 43168 7760 43220 7812
rect 47124 7803 47176 7812
rect 31852 7735 31904 7744
rect 31852 7701 31861 7735
rect 31861 7701 31895 7735
rect 31895 7701 31904 7735
rect 31852 7692 31904 7701
rect 33784 7735 33836 7744
rect 33784 7701 33793 7735
rect 33793 7701 33827 7735
rect 33827 7701 33836 7735
rect 33784 7692 33836 7701
rect 34336 7692 34388 7744
rect 47124 7769 47133 7803
rect 47133 7769 47167 7803
rect 47167 7769 47176 7803
rect 47124 7760 47176 7769
rect 58072 7803 58124 7812
rect 58072 7769 58081 7803
rect 58081 7769 58115 7803
rect 58115 7769 58124 7803
rect 58072 7760 58124 7769
rect 46388 7735 46440 7744
rect 46388 7701 46397 7735
rect 46397 7701 46431 7735
rect 46431 7701 46440 7735
rect 46388 7692 46440 7701
rect 15398 7590 15450 7642
rect 15462 7590 15514 7642
rect 15526 7590 15578 7642
rect 15590 7590 15642 7642
rect 15654 7590 15706 7642
rect 29846 7590 29898 7642
rect 29910 7590 29962 7642
rect 29974 7590 30026 7642
rect 30038 7590 30090 7642
rect 30102 7590 30154 7642
rect 44294 7590 44346 7642
rect 44358 7590 44410 7642
rect 44422 7590 44474 7642
rect 44486 7590 44538 7642
rect 44550 7590 44602 7642
rect 27620 7488 27672 7540
rect 28080 7488 28132 7540
rect 28724 7488 28776 7540
rect 29736 7488 29788 7540
rect 32680 7531 32732 7540
rect 32680 7497 32689 7531
rect 32689 7497 32723 7531
rect 32723 7497 32732 7531
rect 32680 7488 32732 7497
rect 7564 7420 7616 7472
rect 21640 7420 21692 7472
rect 29184 7463 29236 7472
rect 29184 7429 29211 7463
rect 29211 7429 29236 7463
rect 29184 7420 29236 7429
rect 34428 7488 34480 7540
rect 38384 7488 38436 7540
rect 38476 7488 38528 7540
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 28264 7395 28316 7404
rect 28264 7361 28273 7395
rect 28273 7361 28307 7395
rect 28307 7361 28316 7395
rect 28264 7352 28316 7361
rect 28632 7352 28684 7404
rect 29644 7352 29696 7404
rect 27712 7284 27764 7336
rect 28356 7327 28408 7336
rect 27988 7216 28040 7268
rect 28356 7293 28365 7327
rect 28365 7293 28399 7327
rect 28399 7293 28408 7327
rect 28356 7284 28408 7293
rect 28448 7284 28500 7336
rect 30748 7352 30800 7404
rect 39764 7463 39816 7472
rect 39764 7429 39773 7463
rect 39773 7429 39807 7463
rect 39807 7429 39816 7463
rect 39764 7420 39816 7429
rect 31576 7352 31628 7404
rect 33048 7352 33100 7404
rect 34244 7352 34296 7404
rect 37740 7395 37792 7404
rect 31208 7327 31260 7336
rect 31208 7293 31217 7327
rect 31217 7293 31251 7327
rect 31251 7293 31260 7327
rect 31208 7284 31260 7293
rect 31300 7284 31352 7336
rect 34336 7327 34388 7336
rect 34336 7293 34345 7327
rect 34345 7293 34379 7327
rect 34379 7293 34388 7327
rect 34336 7284 34388 7293
rect 33600 7216 33652 7268
rect 36728 7259 36780 7268
rect 36728 7225 36737 7259
rect 36737 7225 36771 7259
rect 36771 7225 36780 7259
rect 37740 7361 37749 7395
rect 37749 7361 37783 7395
rect 37783 7361 37792 7395
rect 37740 7352 37792 7361
rect 40040 7395 40092 7404
rect 40040 7361 40049 7395
rect 40049 7361 40083 7395
rect 40083 7361 40092 7395
rect 41144 7488 41196 7540
rect 44640 7488 44692 7540
rect 44732 7531 44784 7540
rect 44732 7497 44741 7531
rect 44741 7497 44775 7531
rect 44775 7497 44784 7531
rect 44732 7488 44784 7497
rect 46296 7488 46348 7540
rect 46572 7531 46624 7540
rect 46572 7497 46581 7531
rect 46581 7497 46615 7531
rect 46615 7497 46624 7531
rect 46572 7488 46624 7497
rect 40408 7420 40460 7472
rect 41696 7420 41748 7472
rect 43168 7420 43220 7472
rect 45560 7420 45612 7472
rect 47124 7420 47176 7472
rect 40040 7352 40092 7361
rect 41328 7352 41380 7404
rect 42340 7352 42392 7404
rect 45100 7352 45152 7404
rect 45468 7352 45520 7404
rect 45928 7395 45980 7404
rect 45928 7361 45937 7395
rect 45937 7361 45971 7395
rect 45971 7361 45980 7395
rect 45928 7352 45980 7361
rect 38568 7284 38620 7336
rect 39212 7284 39264 7336
rect 45192 7284 45244 7336
rect 36728 7216 36780 7225
rect 28080 7148 28132 7200
rect 29092 7148 29144 7200
rect 29644 7148 29696 7200
rect 34704 7191 34756 7200
rect 34704 7157 34713 7191
rect 34713 7157 34747 7191
rect 34747 7157 34756 7191
rect 34704 7148 34756 7157
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 8302 7046 8354 7098
rect 8366 7046 8418 7098
rect 8430 7046 8482 7098
rect 22622 7046 22674 7098
rect 22686 7046 22738 7098
rect 22750 7046 22802 7098
rect 22814 7046 22866 7098
rect 22878 7046 22930 7098
rect 37070 7046 37122 7098
rect 37134 7046 37186 7098
rect 37198 7046 37250 7098
rect 37262 7046 37314 7098
rect 37326 7046 37378 7098
rect 51518 7046 51570 7098
rect 51582 7046 51634 7098
rect 51646 7046 51698 7098
rect 51710 7046 51762 7098
rect 51774 7046 51826 7098
rect 21640 6987 21692 6996
rect 21640 6953 21649 6987
rect 21649 6953 21683 6987
rect 21683 6953 21692 6987
rect 21640 6944 21692 6953
rect 30472 6944 30524 6996
rect 31208 6944 31260 6996
rect 31852 6944 31904 6996
rect 33784 6944 33836 6996
rect 34704 6944 34756 6996
rect 45100 6987 45152 6996
rect 45100 6953 45109 6987
rect 45109 6953 45143 6987
rect 45143 6953 45152 6987
rect 45100 6944 45152 6953
rect 46388 6944 46440 6996
rect 46480 6987 46532 6996
rect 46480 6953 46489 6987
rect 46489 6953 46523 6987
rect 46523 6953 46532 6987
rect 46480 6944 46532 6953
rect 27988 6919 28040 6928
rect 27988 6885 27997 6919
rect 27997 6885 28031 6919
rect 28031 6885 28040 6919
rect 27988 6876 28040 6885
rect 20536 6808 20588 6860
rect 7932 6740 7984 6792
rect 19524 6740 19576 6792
rect 27620 6808 27672 6860
rect 27804 6740 27856 6792
rect 29460 6808 29512 6860
rect 31576 6808 31628 6860
rect 32220 6851 32272 6860
rect 32220 6817 32229 6851
rect 32229 6817 32263 6851
rect 32263 6817 32272 6851
rect 32220 6808 32272 6817
rect 29092 6740 29144 6792
rect 30196 6740 30248 6792
rect 30472 6783 30524 6792
rect 30472 6749 30481 6783
rect 30481 6749 30515 6783
rect 30515 6749 30524 6783
rect 30472 6740 30524 6749
rect 30564 6783 30616 6792
rect 30564 6749 30573 6783
rect 30573 6749 30607 6783
rect 30607 6749 30616 6783
rect 30840 6783 30892 6792
rect 30564 6740 30616 6749
rect 30840 6749 30849 6783
rect 30849 6749 30883 6783
rect 30883 6749 30892 6783
rect 30840 6740 30892 6749
rect 35072 6876 35124 6928
rect 34244 6808 34296 6860
rect 39028 6851 39080 6860
rect 39028 6817 39037 6851
rect 39037 6817 39071 6851
rect 39071 6817 39080 6851
rect 39028 6808 39080 6817
rect 39856 6808 39908 6860
rect 28356 6715 28408 6724
rect 28356 6681 28365 6715
rect 28365 6681 28399 6715
rect 28399 6681 28408 6715
rect 34428 6740 34480 6792
rect 34520 6740 34572 6792
rect 35072 6740 35124 6792
rect 38476 6740 38528 6792
rect 38844 6740 38896 6792
rect 39120 6783 39172 6792
rect 39120 6749 39129 6783
rect 39129 6749 39163 6783
rect 39163 6749 39172 6783
rect 39120 6740 39172 6749
rect 40408 6783 40460 6792
rect 40408 6749 40417 6783
rect 40417 6749 40451 6783
rect 40451 6749 40460 6783
rect 40408 6740 40460 6749
rect 38016 6715 38068 6724
rect 28356 6672 28408 6681
rect 38016 6681 38025 6715
rect 38025 6681 38059 6715
rect 38059 6681 38068 6715
rect 38016 6672 38068 6681
rect 40684 6672 40736 6724
rect 44088 6740 44140 6792
rect 45560 6740 45612 6792
rect 45928 6740 45980 6792
rect 43076 6672 43128 6724
rect 44732 6672 44784 6724
rect 19708 6647 19760 6656
rect 19708 6613 19717 6647
rect 19717 6613 19751 6647
rect 19751 6613 19760 6647
rect 19708 6604 19760 6613
rect 27712 6604 27764 6656
rect 28264 6647 28316 6656
rect 28264 6613 28273 6647
rect 28273 6613 28307 6647
rect 28307 6613 28316 6647
rect 28264 6604 28316 6613
rect 29184 6604 29236 6656
rect 29368 6604 29420 6656
rect 29736 6647 29788 6656
rect 29736 6613 29745 6647
rect 29745 6613 29779 6647
rect 29779 6613 29788 6647
rect 29736 6604 29788 6613
rect 30656 6647 30708 6656
rect 30656 6613 30665 6647
rect 30665 6613 30699 6647
rect 30699 6613 30708 6647
rect 30656 6604 30708 6613
rect 40408 6604 40460 6656
rect 41880 6647 41932 6656
rect 41880 6613 41889 6647
rect 41889 6613 41923 6647
rect 41923 6613 41932 6647
rect 41880 6604 41932 6613
rect 42892 6604 42944 6656
rect 42984 6604 43036 6656
rect 15398 6502 15450 6554
rect 15462 6502 15514 6554
rect 15526 6502 15578 6554
rect 15590 6502 15642 6554
rect 15654 6502 15706 6554
rect 29846 6502 29898 6554
rect 29910 6502 29962 6554
rect 29974 6502 30026 6554
rect 30038 6502 30090 6554
rect 30102 6502 30154 6554
rect 44294 6502 44346 6554
rect 44358 6502 44410 6554
rect 44422 6502 44474 6554
rect 44486 6502 44538 6554
rect 44550 6502 44602 6554
rect 19524 6443 19576 6452
rect 19524 6409 19533 6443
rect 19533 6409 19567 6443
rect 19567 6409 19576 6443
rect 19524 6400 19576 6409
rect 34428 6400 34480 6452
rect 36728 6443 36780 6452
rect 36728 6409 36737 6443
rect 36737 6409 36771 6443
rect 36771 6409 36780 6443
rect 36728 6400 36780 6409
rect 41880 6400 41932 6452
rect 45928 6400 45980 6452
rect 27804 6332 27856 6384
rect 28264 6332 28316 6384
rect 33600 6375 33652 6384
rect 28080 6264 28132 6316
rect 29368 6307 29420 6316
rect 29368 6273 29377 6307
rect 29377 6273 29411 6307
rect 29411 6273 29420 6307
rect 29368 6264 29420 6273
rect 30472 6264 30524 6316
rect 33600 6341 33609 6375
rect 33609 6341 33643 6375
rect 33643 6341 33652 6375
rect 33600 6332 33652 6341
rect 35900 6332 35952 6384
rect 33232 6264 33284 6316
rect 38200 6332 38252 6384
rect 37924 6307 37976 6316
rect 37924 6273 37933 6307
rect 37933 6273 37967 6307
rect 37967 6273 37976 6307
rect 37924 6264 37976 6273
rect 38752 6307 38804 6316
rect 38752 6273 38761 6307
rect 38761 6273 38795 6307
rect 38795 6273 38804 6307
rect 38752 6264 38804 6273
rect 41788 6332 41840 6384
rect 25964 6196 26016 6248
rect 29460 6196 29512 6248
rect 29736 6196 29788 6248
rect 32404 6196 32456 6248
rect 36636 6196 36688 6248
rect 27712 6128 27764 6180
rect 33232 6128 33284 6180
rect 28724 6060 28776 6112
rect 30196 6060 30248 6112
rect 32220 6060 32272 6112
rect 32588 6060 32640 6112
rect 39856 6264 39908 6316
rect 41512 6264 41564 6316
rect 42892 6264 42944 6316
rect 42984 6307 43036 6316
rect 42984 6273 42993 6307
rect 42993 6273 43027 6307
rect 43027 6273 43036 6307
rect 43996 6307 44048 6316
rect 42984 6264 43036 6273
rect 43996 6273 44005 6307
rect 44005 6273 44039 6307
rect 44039 6273 44048 6307
rect 43996 6264 44048 6273
rect 40684 6196 40736 6248
rect 40592 6128 40644 6180
rect 43628 6171 43680 6180
rect 43628 6137 43637 6171
rect 43637 6137 43671 6171
rect 43671 6137 43680 6171
rect 43628 6128 43680 6137
rect 37740 6060 37792 6112
rect 39028 6103 39080 6112
rect 39028 6069 39037 6103
rect 39037 6069 39071 6103
rect 39071 6069 39080 6103
rect 39028 6060 39080 6069
rect 40132 6060 40184 6112
rect 43076 6060 43128 6112
rect 43536 6060 43588 6112
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 8302 5958 8354 6010
rect 8366 5958 8418 6010
rect 8430 5958 8482 6010
rect 22622 5958 22674 6010
rect 22686 5958 22738 6010
rect 22750 5958 22802 6010
rect 22814 5958 22866 6010
rect 22878 5958 22930 6010
rect 37070 5958 37122 6010
rect 37134 5958 37186 6010
rect 37198 5958 37250 6010
rect 37262 5958 37314 6010
rect 37326 5958 37378 6010
rect 51518 5958 51570 6010
rect 51582 5958 51634 6010
rect 51646 5958 51698 6010
rect 51710 5958 51762 6010
rect 51774 5958 51826 6010
rect 25964 5899 26016 5908
rect 25964 5865 25973 5899
rect 25973 5865 26007 5899
rect 26007 5865 26016 5899
rect 25964 5856 26016 5865
rect 27804 5856 27856 5908
rect 28908 5856 28960 5908
rect 32312 5856 32364 5908
rect 32496 5856 32548 5908
rect 28724 5763 28776 5772
rect 28724 5729 28733 5763
rect 28733 5729 28767 5763
rect 28767 5729 28776 5763
rect 28724 5720 28776 5729
rect 32404 5763 32456 5772
rect 26240 5652 26292 5704
rect 28632 5695 28684 5704
rect 28632 5661 28641 5695
rect 28641 5661 28675 5695
rect 28675 5661 28684 5695
rect 28632 5652 28684 5661
rect 30748 5695 30800 5704
rect 30748 5661 30757 5695
rect 30757 5661 30791 5695
rect 30791 5661 30800 5695
rect 30748 5652 30800 5661
rect 30840 5652 30892 5704
rect 31024 5652 31076 5704
rect 32404 5729 32413 5763
rect 32413 5729 32447 5763
rect 32447 5729 32456 5763
rect 32404 5720 32456 5729
rect 35072 5788 35124 5840
rect 32772 5720 32824 5772
rect 29184 5516 29236 5568
rect 30656 5559 30708 5568
rect 30656 5525 30665 5559
rect 30665 5525 30699 5559
rect 30699 5525 30708 5559
rect 30656 5516 30708 5525
rect 32312 5652 32364 5704
rect 37924 5856 37976 5908
rect 39028 5831 39080 5840
rect 39028 5797 39037 5831
rect 39037 5797 39071 5831
rect 39071 5797 39080 5831
rect 39028 5788 39080 5797
rect 40592 5720 40644 5772
rect 36728 5652 36780 5704
rect 40224 5652 40276 5704
rect 41512 5652 41564 5704
rect 42984 5788 43036 5840
rect 44088 5695 44140 5704
rect 44088 5661 44097 5695
rect 44097 5661 44131 5695
rect 44131 5661 44140 5695
rect 44088 5652 44140 5661
rect 32220 5584 32272 5636
rect 32772 5584 32824 5636
rect 34336 5584 34388 5636
rect 37556 5627 37608 5636
rect 37556 5593 37565 5627
rect 37565 5593 37599 5627
rect 37599 5593 37608 5627
rect 37556 5584 37608 5593
rect 38016 5584 38068 5636
rect 42892 5584 42944 5636
rect 43444 5627 43496 5636
rect 43444 5593 43453 5627
rect 43453 5593 43487 5627
rect 43487 5593 43496 5627
rect 43444 5584 43496 5593
rect 43536 5584 43588 5636
rect 38936 5516 38988 5568
rect 39948 5516 40000 5568
rect 42708 5516 42760 5568
rect 43996 5516 44048 5568
rect 15398 5414 15450 5466
rect 15462 5414 15514 5466
rect 15526 5414 15578 5466
rect 15590 5414 15642 5466
rect 15654 5414 15706 5466
rect 29846 5414 29898 5466
rect 29910 5414 29962 5466
rect 29974 5414 30026 5466
rect 30038 5414 30090 5466
rect 30102 5414 30154 5466
rect 44294 5414 44346 5466
rect 44358 5414 44410 5466
rect 44422 5414 44474 5466
rect 44486 5414 44538 5466
rect 44550 5414 44602 5466
rect 19708 5312 19760 5364
rect 21732 5312 21784 5364
rect 26240 5355 26292 5364
rect 26240 5321 26249 5355
rect 26249 5321 26283 5355
rect 26283 5321 26292 5355
rect 26240 5312 26292 5321
rect 30656 5312 30708 5364
rect 33324 5355 33376 5364
rect 33324 5321 33333 5355
rect 33333 5321 33367 5355
rect 33367 5321 33376 5355
rect 33324 5312 33376 5321
rect 37556 5312 37608 5364
rect 40040 5312 40092 5364
rect 40316 5355 40368 5364
rect 40316 5321 40325 5355
rect 40325 5321 40359 5355
rect 40359 5321 40368 5355
rect 40316 5312 40368 5321
rect 41512 5312 41564 5364
rect 30288 5244 30340 5296
rect 34336 5244 34388 5296
rect 35808 5244 35860 5296
rect 38936 5244 38988 5296
rect 41604 5287 41656 5296
rect 41604 5253 41613 5287
rect 41613 5253 41647 5287
rect 41647 5253 41656 5287
rect 41604 5244 41656 5253
rect 41788 5287 41840 5296
rect 41788 5253 41797 5287
rect 41797 5253 41831 5287
rect 41831 5253 41840 5287
rect 41788 5244 41840 5253
rect 25872 5219 25924 5228
rect 25872 5185 25881 5219
rect 25881 5185 25915 5219
rect 25915 5185 25924 5219
rect 25872 5176 25924 5185
rect 26976 5176 27028 5228
rect 29184 5108 29236 5160
rect 29644 5176 29696 5228
rect 30472 5176 30524 5228
rect 31024 5219 31076 5228
rect 31024 5185 31033 5219
rect 31033 5185 31067 5219
rect 31067 5185 31076 5219
rect 31024 5176 31076 5185
rect 32312 5219 32364 5228
rect 32312 5185 32321 5219
rect 32321 5185 32355 5219
rect 32355 5185 32364 5219
rect 32312 5176 32364 5185
rect 32496 5219 32548 5228
rect 32496 5185 32505 5219
rect 32505 5185 32539 5219
rect 32539 5185 32548 5219
rect 32496 5176 32548 5185
rect 32588 5219 32640 5228
rect 32588 5185 32597 5219
rect 32597 5185 32631 5219
rect 32631 5185 32640 5219
rect 37648 5219 37700 5228
rect 32588 5176 32640 5185
rect 37648 5185 37657 5219
rect 37657 5185 37691 5219
rect 37691 5185 37700 5219
rect 37648 5176 37700 5185
rect 38108 5176 38160 5228
rect 40224 5176 40276 5228
rect 41512 5219 41564 5228
rect 41512 5185 41521 5219
rect 41521 5185 41555 5219
rect 41555 5185 41564 5219
rect 41512 5176 41564 5185
rect 43076 5176 43128 5228
rect 30380 5108 30432 5160
rect 30564 5108 30616 5160
rect 31484 5108 31536 5160
rect 32036 5108 32088 5160
rect 24768 5040 24820 5092
rect 33048 5040 33100 5092
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 24860 4972 24912 5024
rect 32128 5015 32180 5024
rect 32128 4981 32137 5015
rect 32137 4981 32171 5015
rect 32171 4981 32180 5015
rect 32128 4972 32180 4981
rect 33232 5108 33284 5160
rect 35072 5151 35124 5160
rect 35072 5117 35081 5151
rect 35081 5117 35115 5151
rect 35115 5117 35124 5151
rect 35072 5108 35124 5117
rect 37740 5151 37792 5160
rect 37740 5117 37749 5151
rect 37749 5117 37783 5151
rect 37783 5117 37792 5151
rect 37740 5108 37792 5117
rect 38292 5151 38344 5160
rect 38292 5117 38301 5151
rect 38301 5117 38335 5151
rect 38335 5117 38344 5151
rect 38292 5108 38344 5117
rect 43444 5108 43496 5160
rect 35256 5040 35308 5092
rect 39856 5040 39908 5092
rect 36636 4972 36688 5024
rect 37556 4972 37608 5024
rect 39948 4972 40000 5024
rect 43536 4972 43588 5024
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 8302 4870 8354 4922
rect 8366 4870 8418 4922
rect 8430 4870 8482 4922
rect 22622 4870 22674 4922
rect 22686 4870 22738 4922
rect 22750 4870 22802 4922
rect 22814 4870 22866 4922
rect 22878 4870 22930 4922
rect 37070 4870 37122 4922
rect 37134 4870 37186 4922
rect 37198 4870 37250 4922
rect 37262 4870 37314 4922
rect 37326 4870 37378 4922
rect 51518 4870 51570 4922
rect 51582 4870 51634 4922
rect 51646 4870 51698 4922
rect 51710 4870 51762 4922
rect 51774 4870 51826 4922
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 25872 4811 25924 4820
rect 25872 4777 25881 4811
rect 25881 4777 25915 4811
rect 25915 4777 25924 4811
rect 25872 4768 25924 4777
rect 26332 4700 26384 4752
rect 24860 4607 24912 4616
rect 24860 4573 24869 4607
rect 24869 4573 24903 4607
rect 24903 4573 24912 4607
rect 24860 4564 24912 4573
rect 29644 4632 29696 4684
rect 29184 4564 29236 4616
rect 25412 4539 25464 4548
rect 25412 4505 25421 4539
rect 25421 4505 25455 4539
rect 25455 4505 25464 4539
rect 25412 4496 25464 4505
rect 26332 4539 26384 4548
rect 26332 4505 26341 4539
rect 26341 4505 26375 4539
rect 26375 4505 26384 4539
rect 26332 4496 26384 4505
rect 32496 4768 32548 4820
rect 33140 4768 33192 4820
rect 37648 4768 37700 4820
rect 39948 4811 40000 4820
rect 31392 4632 31444 4684
rect 31484 4564 31536 4616
rect 32036 4607 32088 4616
rect 32036 4573 32045 4607
rect 32045 4573 32079 4607
rect 32079 4573 32088 4607
rect 32036 4564 32088 4573
rect 33140 4632 33192 4684
rect 38200 4675 38252 4684
rect 38200 4641 38209 4675
rect 38209 4641 38243 4675
rect 38243 4641 38252 4675
rect 38200 4632 38252 4641
rect 39948 4777 39957 4811
rect 39957 4777 39991 4811
rect 39991 4777 40000 4811
rect 39948 4768 40000 4777
rect 41512 4768 41564 4820
rect 41604 4700 41656 4752
rect 39028 4632 39080 4684
rect 42432 4632 42484 4684
rect 27160 4428 27212 4480
rect 27252 4428 27304 4480
rect 29644 4471 29696 4480
rect 29644 4437 29653 4471
rect 29653 4437 29687 4471
rect 29687 4437 29696 4471
rect 29644 4428 29696 4437
rect 31760 4496 31812 4548
rect 35256 4539 35308 4548
rect 35256 4505 35265 4539
rect 35265 4505 35299 4539
rect 35299 4505 35308 4539
rect 35256 4496 35308 4505
rect 38108 4564 38160 4616
rect 37740 4539 37792 4548
rect 37740 4505 37749 4539
rect 37749 4505 37783 4539
rect 37783 4505 37792 4539
rect 38752 4564 38804 4616
rect 39856 4564 39908 4616
rect 37740 4496 37792 4505
rect 41328 4496 41380 4548
rect 43628 4496 43680 4548
rect 15398 4326 15450 4378
rect 15462 4326 15514 4378
rect 15526 4326 15578 4378
rect 15590 4326 15642 4378
rect 15654 4326 15706 4378
rect 29846 4326 29898 4378
rect 29910 4326 29962 4378
rect 29974 4326 30026 4378
rect 30038 4326 30090 4378
rect 30102 4326 30154 4378
rect 44294 4326 44346 4378
rect 44358 4326 44410 4378
rect 44422 4326 44474 4378
rect 44486 4326 44538 4378
rect 44550 4326 44602 4378
rect 26976 4267 27028 4276
rect 26976 4233 26985 4267
rect 26985 4233 27019 4267
rect 27019 4233 27028 4267
rect 26976 4224 27028 4233
rect 31760 4224 31812 4276
rect 34428 4224 34480 4276
rect 27252 4156 27304 4208
rect 35256 4224 35308 4276
rect 40592 4267 40644 4276
rect 40592 4233 40601 4267
rect 40601 4233 40635 4267
rect 40635 4233 40644 4267
rect 40592 4224 40644 4233
rect 13636 4088 13688 4140
rect 14280 4088 14332 4140
rect 27160 4131 27212 4140
rect 27160 4097 27169 4131
rect 27169 4097 27203 4131
rect 27203 4097 27212 4131
rect 27160 4088 27212 4097
rect 25320 4020 25372 4072
rect 25412 3952 25464 4004
rect 23112 3927 23164 3936
rect 23112 3893 23121 3927
rect 23121 3893 23155 3927
rect 23155 3893 23164 3927
rect 23112 3884 23164 3893
rect 25320 3927 25372 3936
rect 25320 3893 25329 3927
rect 25329 3893 25363 3927
rect 25363 3893 25372 3927
rect 25320 3884 25372 3893
rect 29184 3927 29236 3936
rect 29184 3893 29193 3927
rect 29193 3893 29227 3927
rect 29227 3893 29236 3927
rect 29184 3884 29236 3893
rect 32128 4088 32180 4140
rect 32404 4088 32456 4140
rect 37740 4088 37792 4140
rect 40408 4156 40460 4208
rect 41328 4156 41380 4208
rect 42432 4131 42484 4140
rect 34888 4063 34940 4072
rect 34888 4029 34897 4063
rect 34897 4029 34931 4063
rect 34931 4029 34940 4063
rect 34888 4020 34940 4029
rect 34520 3952 34572 4004
rect 36636 4063 36688 4072
rect 36636 4029 36645 4063
rect 36645 4029 36679 4063
rect 36679 4029 36688 4063
rect 36636 4020 36688 4029
rect 37556 4063 37608 4072
rect 37556 4029 37565 4063
rect 37565 4029 37599 4063
rect 37599 4029 37608 4063
rect 37556 4020 37608 4029
rect 40316 4020 40368 4072
rect 42432 4097 42441 4131
rect 42441 4097 42475 4131
rect 42475 4097 42484 4131
rect 42432 4088 42484 4097
rect 48688 4131 48740 4140
rect 48688 4097 48697 4131
rect 48697 4097 48731 4131
rect 48731 4097 48740 4131
rect 48688 4088 48740 4097
rect 42708 4063 42760 4072
rect 42708 4029 42717 4063
rect 42717 4029 42751 4063
rect 42751 4029 42760 4063
rect 42708 4020 42760 4029
rect 43076 4020 43128 4072
rect 31944 3884 31996 3936
rect 32588 3884 32640 3936
rect 34428 3927 34480 3936
rect 34428 3893 34437 3927
rect 34437 3893 34471 3927
rect 34471 3893 34480 3927
rect 48872 3927 48924 3936
rect 34428 3884 34480 3893
rect 48872 3893 48881 3927
rect 48881 3893 48915 3927
rect 48915 3893 48924 3927
rect 48872 3884 48924 3893
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 8302 3782 8354 3834
rect 8366 3782 8418 3834
rect 8430 3782 8482 3834
rect 22622 3782 22674 3834
rect 22686 3782 22738 3834
rect 22750 3782 22802 3834
rect 22814 3782 22866 3834
rect 22878 3782 22930 3834
rect 37070 3782 37122 3834
rect 37134 3782 37186 3834
rect 37198 3782 37250 3834
rect 37262 3782 37314 3834
rect 37326 3782 37378 3834
rect 51518 3782 51570 3834
rect 51582 3782 51634 3834
rect 51646 3782 51698 3834
rect 51710 3782 51762 3834
rect 51774 3782 51826 3834
rect 26332 3680 26384 3732
rect 23112 3544 23164 3596
rect 25320 3476 25372 3528
rect 27252 3408 27304 3460
rect 29184 3680 29236 3732
rect 32588 3680 32640 3732
rect 34428 3680 34480 3732
rect 30380 3612 30432 3664
rect 28080 3544 28132 3596
rect 48688 3680 48740 3732
rect 35072 3612 35124 3664
rect 41788 3612 41840 3664
rect 40224 3544 40276 3596
rect 35164 3408 35216 3460
rect 40132 3451 40184 3460
rect 33048 3340 33100 3392
rect 40132 3417 40141 3451
rect 40141 3417 40175 3451
rect 40175 3417 40184 3451
rect 40132 3408 40184 3417
rect 40408 3408 40460 3460
rect 15398 3238 15450 3290
rect 15462 3238 15514 3290
rect 15526 3238 15578 3290
rect 15590 3238 15642 3290
rect 15654 3238 15706 3290
rect 29846 3238 29898 3290
rect 29910 3238 29962 3290
rect 29974 3238 30026 3290
rect 30038 3238 30090 3290
rect 30102 3238 30154 3290
rect 44294 3238 44346 3290
rect 44358 3238 44410 3290
rect 44422 3238 44474 3290
rect 44486 3238 44538 3290
rect 44550 3238 44602 3290
rect 14280 3136 14332 3188
rect 29644 3136 29696 3188
rect 44180 3136 44232 3188
rect 38016 3068 38068 3120
rect 41236 3068 41288 3120
rect 19708 3000 19760 3052
rect 27896 3043 27948 3052
rect 27896 3009 27905 3043
rect 27905 3009 27939 3043
rect 27939 3009 27948 3043
rect 27896 3000 27948 3009
rect 32404 3000 32456 3052
rect 34888 3000 34940 3052
rect 48872 3000 48924 3052
rect 29184 2932 29236 2984
rect 29552 2864 29604 2916
rect 19708 2796 19760 2848
rect 33784 2796 33836 2848
rect 53104 2864 53156 2916
rect 52828 2796 52880 2848
rect 58072 2839 58124 2848
rect 58072 2805 58081 2839
rect 58081 2805 58115 2839
rect 58115 2805 58124 2839
rect 58072 2796 58124 2805
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 8302 2694 8354 2746
rect 8366 2694 8418 2746
rect 8430 2694 8482 2746
rect 22622 2694 22674 2746
rect 22686 2694 22738 2746
rect 22750 2694 22802 2746
rect 22814 2694 22866 2746
rect 22878 2694 22930 2746
rect 37070 2694 37122 2746
rect 37134 2694 37186 2746
rect 37198 2694 37250 2746
rect 37262 2694 37314 2746
rect 37326 2694 37378 2746
rect 51518 2694 51570 2746
rect 51582 2694 51634 2746
rect 51646 2694 51698 2746
rect 51710 2694 51762 2746
rect 51774 2694 51826 2746
rect 37832 2592 37884 2644
rect 13820 2524 13872 2576
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 4528 2388 4580 2440
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 14280 2388 14332 2397
rect 19708 2431 19760 2440
rect 19708 2397 19717 2431
rect 19717 2397 19751 2431
rect 19751 2397 19760 2431
rect 19708 2388 19760 2397
rect 29552 2431 29604 2440
rect 9680 2320 9732 2372
rect 20 2252 72 2304
rect 16304 2320 16356 2372
rect 29552 2397 29561 2431
rect 29561 2397 29595 2431
rect 29595 2397 29604 2431
rect 29552 2388 29604 2397
rect 33784 2431 33836 2440
rect 33784 2397 33793 2431
rect 33793 2397 33827 2431
rect 33827 2397 33836 2431
rect 33784 2388 33836 2397
rect 41236 2592 41288 2644
rect 53104 2567 53156 2576
rect 53104 2533 53113 2567
rect 53113 2533 53147 2567
rect 53147 2533 53156 2567
rect 53104 2524 53156 2533
rect 43168 2388 43220 2440
rect 48412 2431 48464 2440
rect 48412 2397 48421 2431
rect 48421 2397 48455 2431
rect 48455 2397 48464 2431
rect 48412 2388 48464 2397
rect 57888 2431 57940 2440
rect 57888 2397 57897 2431
rect 57897 2397 57931 2431
rect 57931 2397 57940 2431
rect 57888 2388 57940 2397
rect 41420 2320 41472 2372
rect 52828 2320 52880 2372
rect 14188 2252 14240 2304
rect 19340 2252 19392 2304
rect 23848 2252 23900 2304
rect 29000 2252 29052 2304
rect 33508 2252 33560 2304
rect 38660 2252 38712 2304
rect 48320 2252 48372 2304
rect 57980 2252 58032 2304
rect 15398 2150 15450 2202
rect 15462 2150 15514 2202
rect 15526 2150 15578 2202
rect 15590 2150 15642 2202
rect 15654 2150 15706 2202
rect 29846 2150 29898 2202
rect 29910 2150 29962 2202
rect 29974 2150 30026 2202
rect 30038 2150 30090 2202
rect 30102 2150 30154 2202
rect 44294 2150 44346 2202
rect 44358 2150 44410 2202
rect 44422 2150 44474 2202
rect 44486 2150 44538 2202
rect 44550 2150 44602 2202
<< metal2 >>
rect 1490 35456 1546 35465
rect 1490 35391 1546 35400
rect 1504 33658 1532 35391
rect 4526 35306 4582 36000
rect 4526 35278 4844 35306
rect 4526 35200 4582 35278
rect 4816 33658 4844 35278
rect 9034 35200 9090 36000
rect 14186 35306 14242 36000
rect 14186 35278 14412 35306
rect 14186 35200 14242 35278
rect 9048 33658 9076 35200
rect 14384 33658 14412 35278
rect 18694 35200 18750 36000
rect 23846 35200 23902 36000
rect 28354 35306 28410 36000
rect 33506 35306 33562 36000
rect 28354 35278 28580 35306
rect 28354 35200 28410 35278
rect 15398 33756 15706 33765
rect 15398 33754 15404 33756
rect 15460 33754 15484 33756
rect 15540 33754 15564 33756
rect 15620 33754 15644 33756
rect 15700 33754 15706 33756
rect 15460 33702 15462 33754
rect 15642 33702 15644 33754
rect 15398 33700 15404 33702
rect 15460 33700 15484 33702
rect 15540 33700 15564 33702
rect 15620 33700 15644 33702
rect 15700 33700 15706 33702
rect 15398 33691 15706 33700
rect 18708 33658 18736 35200
rect 1492 33652 1544 33658
rect 1492 33594 1544 33600
rect 4804 33652 4856 33658
rect 4804 33594 4856 33600
rect 9036 33652 9088 33658
rect 9036 33594 9088 33600
rect 14372 33652 14424 33658
rect 14372 33594 14424 33600
rect 18696 33652 18748 33658
rect 18696 33594 18748 33600
rect 23860 33522 23888 35200
rect 28552 33590 28580 35278
rect 33506 35278 33824 35306
rect 33506 35200 33562 35278
rect 29846 33756 30154 33765
rect 29846 33754 29852 33756
rect 29908 33754 29932 33756
rect 29988 33754 30012 33756
rect 30068 33754 30092 33756
rect 30148 33754 30154 33756
rect 29908 33702 29910 33754
rect 30090 33702 30092 33754
rect 29846 33700 29852 33702
rect 29908 33700 29932 33702
rect 29988 33700 30012 33702
rect 30068 33700 30092 33702
rect 30148 33700 30154 33702
rect 29846 33691 30154 33700
rect 33796 33658 33824 35278
rect 38658 35200 38714 36000
rect 43166 35306 43222 36000
rect 48318 35306 48374 36000
rect 52826 35306 52882 36000
rect 43166 35278 43300 35306
rect 43166 35200 43222 35278
rect 38672 33658 38700 35200
rect 43272 33658 43300 35278
rect 48318 35278 48636 35306
rect 48318 35200 48374 35278
rect 44294 33756 44602 33765
rect 44294 33754 44300 33756
rect 44356 33754 44380 33756
rect 44436 33754 44460 33756
rect 44516 33754 44540 33756
rect 44596 33754 44602 33756
rect 44356 33702 44358 33754
rect 44538 33702 44540 33754
rect 44294 33700 44300 33702
rect 44356 33700 44380 33702
rect 44436 33700 44460 33702
rect 44516 33700 44540 33702
rect 44596 33700 44602 33702
rect 44294 33691 44602 33700
rect 48608 33658 48636 35278
rect 52826 35278 53144 35306
rect 52826 35200 52882 35278
rect 53116 33658 53144 35278
rect 57978 35200 58034 36000
rect 33784 33652 33836 33658
rect 33784 33594 33836 33600
rect 38660 33652 38712 33658
rect 38660 33594 38712 33600
rect 43260 33652 43312 33658
rect 43260 33594 43312 33600
rect 48596 33652 48648 33658
rect 48596 33594 48648 33600
rect 53104 33652 53156 33658
rect 53104 33594 53156 33600
rect 28540 33584 28592 33590
rect 57992 33538 58020 35200
rect 28540 33526 28592 33532
rect 57808 33522 58020 33538
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 4620 33516 4672 33522
rect 4620 33458 4672 33464
rect 9404 33516 9456 33522
rect 9404 33458 9456 33464
rect 17224 33516 17276 33522
rect 17224 33458 17276 33464
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 33600 33516 33652 33522
rect 33600 33458 33652 33464
rect 38936 33516 38988 33522
rect 38936 33458 38988 33464
rect 43904 33516 43956 33522
rect 43904 33458 43956 33464
rect 48412 33516 48464 33522
rect 48412 33458 48464 33464
rect 52644 33516 52696 33522
rect 52644 33458 52696 33464
rect 57796 33516 58020 33522
rect 57848 33510 58020 33516
rect 57796 33458 57848 33464
rect 1688 30938 1716 33458
rect 4632 33114 4660 33458
rect 6828 33312 6880 33318
rect 6828 33254 6880 33260
rect 8024 33312 8076 33318
rect 8024 33254 8076 33260
rect 6840 33130 6868 33254
rect 4620 33108 4672 33114
rect 6840 33102 6960 33130
rect 4620 33050 4672 33056
rect 4436 32904 4488 32910
rect 4436 32846 4488 32852
rect 5172 32904 5224 32910
rect 5172 32846 5224 32852
rect 5448 32904 5500 32910
rect 5448 32846 5500 32852
rect 6552 32904 6604 32910
rect 6552 32846 6604 32852
rect 2780 32428 2832 32434
rect 2780 32370 2832 32376
rect 1768 32360 1820 32366
rect 1768 32302 1820 32308
rect 1780 31822 1808 32302
rect 1768 31816 1820 31822
rect 1768 31758 1820 31764
rect 1676 30932 1728 30938
rect 1676 30874 1728 30880
rect 1490 30696 1546 30705
rect 1490 30631 1546 30640
rect 1504 30598 1532 30631
rect 1492 30592 1544 30598
rect 1492 30534 1544 30540
rect 2504 29708 2556 29714
rect 2504 29650 2556 29656
rect 2516 29170 2544 29650
rect 2792 29238 2820 32370
rect 4448 32230 4476 32846
rect 3056 32224 3108 32230
rect 3056 32166 3108 32172
rect 4436 32224 4488 32230
rect 4436 32166 4488 32172
rect 3068 31414 3096 32166
rect 3056 31408 3108 31414
rect 3056 31350 3108 31356
rect 3068 30734 3096 31350
rect 2872 30728 2924 30734
rect 2872 30670 2924 30676
rect 3056 30728 3108 30734
rect 3056 30670 3108 30676
rect 2780 29232 2832 29238
rect 2780 29174 2832 29180
rect 2504 29164 2556 29170
rect 2504 29106 2556 29112
rect 2320 28960 2372 28966
rect 2320 28902 2372 28908
rect 2332 28218 2360 28902
rect 2320 28212 2372 28218
rect 2320 28154 2372 28160
rect 2516 28014 2544 29106
rect 2792 28150 2820 29174
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 1860 28008 1912 28014
rect 1860 27950 1912 27956
rect 2504 28008 2556 28014
rect 2504 27950 2556 27956
rect 1676 26240 1728 26246
rect 1676 26182 1728 26188
rect 1688 25974 1716 26182
rect 1676 25968 1728 25974
rect 1676 25910 1728 25916
rect 1490 25256 1546 25265
rect 1490 25191 1546 25200
rect 1504 25158 1532 25191
rect 1492 25152 1544 25158
rect 1492 25094 1544 25100
rect 1872 10810 1900 27950
rect 2884 27538 2912 30670
rect 4160 30048 4212 30054
rect 4160 29990 4212 29996
rect 4068 29572 4120 29578
rect 4068 29514 4120 29520
rect 3240 29504 3292 29510
rect 3240 29446 3292 29452
rect 3252 29238 3280 29446
rect 4080 29306 4108 29514
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 4172 29238 4200 29990
rect 3240 29232 3292 29238
rect 3240 29174 3292 29180
rect 4160 29232 4212 29238
rect 4160 29174 4212 29180
rect 2872 27532 2924 27538
rect 2872 27474 2924 27480
rect 2504 27396 2556 27402
rect 2504 27338 2556 27344
rect 3884 27396 3936 27402
rect 3884 27338 3936 27344
rect 2516 27130 2544 27338
rect 3700 27328 3752 27334
rect 3700 27270 3752 27276
rect 2504 27124 2556 27130
rect 2504 27066 2556 27072
rect 2412 26784 2464 26790
rect 2412 26726 2464 26732
rect 2424 25294 2452 26726
rect 2872 26376 2924 26382
rect 2872 26318 2924 26324
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 2412 25288 2464 25294
rect 2412 25230 2464 25236
rect 2424 24857 2452 25230
rect 2410 24848 2466 24857
rect 2410 24783 2466 24792
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 2228 24608 2280 24614
rect 2228 24550 2280 24556
rect 1964 23202 1992 24550
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 2056 23730 2084 24006
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 2240 23526 2268 24550
rect 2792 24070 2820 25842
rect 2884 25770 2912 26318
rect 3056 26240 3108 26246
rect 3056 26182 3108 26188
rect 2872 25764 2924 25770
rect 2872 25706 2924 25712
rect 3068 25702 3096 26182
rect 3712 25906 3740 27270
rect 3896 27062 3924 27338
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 27062 4108 27270
rect 4172 27130 4200 29174
rect 4344 28484 4396 28490
rect 4344 28426 4396 28432
rect 4252 28144 4304 28150
rect 4252 28086 4304 28092
rect 4264 27985 4292 28086
rect 4250 27976 4306 27985
rect 4250 27911 4306 27920
rect 4264 27606 4292 27911
rect 4356 27878 4384 28426
rect 4344 27872 4396 27878
rect 4344 27814 4396 27820
rect 4252 27600 4304 27606
rect 4252 27542 4304 27548
rect 4252 27464 4304 27470
rect 4356 27418 4384 27814
rect 4304 27412 4384 27418
rect 4252 27406 4384 27412
rect 4264 27390 4384 27406
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 3884 27056 3936 27062
rect 3884 26998 3936 27004
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3804 26586 3832 26930
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 4080 26450 4108 26794
rect 4068 26444 4120 26450
rect 4068 26386 4120 26392
rect 4080 26234 4108 26386
rect 4264 26234 4292 27390
rect 4448 26790 4476 32166
rect 5184 31822 5212 32846
rect 5460 32502 5488 32846
rect 6368 32768 6420 32774
rect 6368 32710 6420 32716
rect 5448 32496 5500 32502
rect 5448 32438 5500 32444
rect 5460 31822 5488 32438
rect 5172 31816 5224 31822
rect 5172 31758 5224 31764
rect 5448 31816 5500 31822
rect 5448 31758 5500 31764
rect 6184 31816 6236 31822
rect 6184 31758 6236 31764
rect 4620 31680 4672 31686
rect 4620 31622 4672 31628
rect 4632 31142 4660 31622
rect 5460 31346 5488 31758
rect 5816 31408 5868 31414
rect 5816 31350 5868 31356
rect 5448 31340 5500 31346
rect 5448 31282 5500 31288
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4632 30734 4660 31078
rect 5460 30734 5488 31282
rect 5828 30938 5856 31350
rect 6196 31346 6224 31758
rect 6380 31686 6408 32710
rect 6564 32570 6592 32846
rect 6932 32842 6960 33102
rect 6920 32836 6972 32842
rect 6920 32778 6972 32784
rect 7012 32768 7064 32774
rect 6932 32716 7012 32722
rect 6932 32710 7064 32716
rect 6932 32694 7052 32710
rect 6552 32564 6604 32570
rect 6552 32506 6604 32512
rect 6564 31822 6592 32506
rect 6932 32366 6960 32694
rect 7012 32496 7064 32502
rect 7012 32438 7064 32444
rect 7932 32496 7984 32502
rect 7932 32438 7984 32444
rect 6920 32360 6972 32366
rect 6920 32302 6972 32308
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6368 31680 6420 31686
rect 6368 31622 6420 31628
rect 6380 31414 6408 31622
rect 6368 31408 6420 31414
rect 6368 31350 6420 31356
rect 6184 31340 6236 31346
rect 6184 31282 6236 31288
rect 5816 30932 5868 30938
rect 5816 30874 5868 30880
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 5448 30728 5500 30734
rect 5448 30670 5500 30676
rect 4632 30598 4660 30670
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4632 30190 4660 30534
rect 5460 30258 5488 30670
rect 5828 30394 5856 30874
rect 6196 30734 6224 31282
rect 6564 30734 6592 31758
rect 6828 30932 6880 30938
rect 6828 30874 6880 30880
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 6196 30394 6224 30670
rect 5816 30388 5868 30394
rect 5816 30330 5868 30336
rect 6184 30388 6236 30394
rect 6184 30330 6236 30336
rect 6564 30258 6592 30670
rect 6840 30258 6868 30874
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 6552 30252 6604 30258
rect 6552 30194 6604 30200
rect 6828 30252 6880 30258
rect 6828 30194 6880 30200
rect 4620 30184 4672 30190
rect 4620 30126 4672 30132
rect 6932 29782 6960 32302
rect 7024 30326 7052 32438
rect 7656 31680 7708 31686
rect 7656 31622 7708 31628
rect 7668 31346 7696 31622
rect 7656 31340 7708 31346
rect 7656 31282 7708 31288
rect 7668 31142 7696 31282
rect 7656 31136 7708 31142
rect 7656 31078 7708 31084
rect 7668 30598 7696 31078
rect 7656 30592 7708 30598
rect 7656 30534 7708 30540
rect 7012 30320 7064 30326
rect 7012 30262 7064 30268
rect 6920 29776 6972 29782
rect 6920 29718 6972 29724
rect 6000 29640 6052 29646
rect 6000 29582 6052 29588
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 5368 29034 5396 29446
rect 5356 29028 5408 29034
rect 5356 28970 5408 28976
rect 4988 28960 5040 28966
rect 4988 28902 5040 28908
rect 5000 28694 5028 28902
rect 4988 28688 5040 28694
rect 4988 28630 5040 28636
rect 5368 28558 5396 28970
rect 6012 28762 6040 29582
rect 7024 29578 7052 30262
rect 7668 30054 7696 30534
rect 7840 30252 7892 30258
rect 7840 30194 7892 30200
rect 7656 30048 7708 30054
rect 7656 29990 7708 29996
rect 7012 29572 7064 29578
rect 7012 29514 7064 29520
rect 6276 29504 6328 29510
rect 6276 29446 6328 29452
rect 6184 29028 6236 29034
rect 6184 28970 6236 28976
rect 6000 28756 6052 28762
rect 6000 28698 6052 28704
rect 6196 28558 6224 28970
rect 6288 28558 6316 29446
rect 7024 29306 7052 29514
rect 7012 29300 7064 29306
rect 7012 29242 7064 29248
rect 6736 29232 6788 29238
rect 6736 29174 6788 29180
rect 7024 29186 7052 29242
rect 6368 28960 6420 28966
rect 6368 28902 6420 28908
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 6276 28552 6328 28558
rect 6276 28494 6328 28500
rect 6288 28150 6316 28494
rect 6380 28218 6408 28902
rect 6748 28558 6776 29174
rect 7024 29158 7144 29186
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 7024 28558 7052 29038
rect 6736 28552 6788 28558
rect 6736 28494 6788 28500
rect 7012 28552 7064 28558
rect 7012 28494 7064 28500
rect 6460 28416 6512 28422
rect 6460 28358 6512 28364
rect 6472 28218 6500 28358
rect 6368 28212 6420 28218
rect 6368 28154 6420 28160
rect 6460 28212 6512 28218
rect 6460 28154 6512 28160
rect 6276 28144 6328 28150
rect 6276 28086 6328 28092
rect 7116 28082 7144 29158
rect 7668 28490 7696 29990
rect 7852 28762 7880 30194
rect 7840 28756 7892 28762
rect 7840 28698 7892 28704
rect 7656 28484 7708 28490
rect 7656 28426 7708 28432
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 7104 28076 7156 28082
rect 7104 28018 7156 28024
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5460 27130 5488 27406
rect 5552 27130 5580 28018
rect 6644 28008 6696 28014
rect 6644 27950 6696 27956
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 4436 26784 4488 26790
rect 4436 26726 4488 26732
rect 5552 26450 5580 27066
rect 5908 26512 5960 26518
rect 5908 26454 5960 26460
rect 5540 26444 5592 26450
rect 5540 26386 5592 26392
rect 5724 26444 5776 26450
rect 5724 26386 5776 26392
rect 5264 26308 5316 26314
rect 5264 26250 5316 26256
rect 3988 26206 4108 26234
rect 4172 26206 4292 26234
rect 3988 26042 4016 26206
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 3608 25696 3660 25702
rect 3608 25638 3660 25644
rect 3976 25696 4028 25702
rect 3976 25638 4028 25644
rect 3068 25140 3096 25638
rect 3148 25152 3200 25158
rect 3068 25112 3148 25140
rect 3148 25094 3200 25100
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3056 24676 3108 24682
rect 3056 24618 3108 24624
rect 2872 24132 2924 24138
rect 2872 24074 2924 24080
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2228 23520 2280 23526
rect 2228 23462 2280 23468
rect 2042 23216 2098 23225
rect 1964 23174 2042 23202
rect 2042 23151 2098 23160
rect 2056 23118 2084 23151
rect 2240 23118 2268 23462
rect 2884 23254 2912 24074
rect 2964 23792 3016 23798
rect 2964 23734 3016 23740
rect 2872 23248 2924 23254
rect 2872 23190 2924 23196
rect 2044 23112 2096 23118
rect 2044 23054 2096 23060
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2240 22098 2268 23054
rect 2780 22976 2832 22982
rect 2976 22930 3004 23734
rect 3068 23730 3096 24618
rect 3160 24206 3188 25094
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 2780 22918 2832 22924
rect 2228 22092 2280 22098
rect 2228 22034 2280 22040
rect 2792 20466 2820 22918
rect 2884 22902 3004 22930
rect 2884 22030 2912 22902
rect 3068 22794 3096 23666
rect 2976 22766 3096 22794
rect 2976 22506 3004 22766
rect 3056 22704 3108 22710
rect 3056 22646 3108 22652
rect 2964 22500 3016 22506
rect 2964 22442 3016 22448
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2884 21622 2912 21830
rect 2872 21616 2924 21622
rect 2872 21558 2924 21564
rect 2976 21146 3004 22442
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2976 20505 3004 20538
rect 2962 20496 3018 20505
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2780 20460 2832 20466
rect 2962 20431 3018 20440
rect 2780 20402 2832 20408
rect 2148 19854 2176 20402
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 2148 19378 2176 19790
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 2148 18766 2176 19314
rect 2240 19310 2268 19858
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 18834 2268 19246
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2148 18290 2176 18702
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2148 17882 2176 18226
rect 2240 18222 2268 18770
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 2884 17746 2912 20334
rect 3068 18766 3096 22646
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 3068 17678 3096 18702
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17270 1992 17478
rect 1952 17264 2004 17270
rect 1952 17206 2004 17212
rect 3068 17066 3096 17614
rect 3056 17060 3108 17066
rect 3056 17002 3108 17008
rect 3160 16998 3188 24142
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3344 23730 3372 24074
rect 3528 24070 3556 25094
rect 3620 24750 3648 25638
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3332 23724 3384 23730
rect 3332 23666 3384 23672
rect 3240 23588 3292 23594
rect 3240 23530 3292 23536
rect 3252 23186 3280 23530
rect 3240 23180 3292 23186
rect 3240 23122 3292 23128
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 3252 21010 3280 21966
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 3240 21004 3292 21010
rect 3240 20946 3292 20952
rect 3148 16992 3200 16998
rect 3148 16934 3200 16940
rect 3344 16182 3372 21422
rect 3528 17270 3556 24006
rect 3712 21894 3740 24754
rect 3792 24064 3844 24070
rect 3792 24006 3844 24012
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3620 21146 3648 21422
rect 3608 21140 3660 21146
rect 3608 21082 3660 21088
rect 3620 20602 3648 21082
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3712 19854 3740 21830
rect 3804 20398 3832 24006
rect 3988 23730 4016 25638
rect 4172 24274 4200 26206
rect 5276 25906 5304 26250
rect 5264 25900 5316 25906
rect 5264 25842 5316 25848
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 4804 25764 4856 25770
rect 4804 25706 4856 25712
rect 4344 25220 4396 25226
rect 4344 25162 4396 25168
rect 4356 24954 4384 25162
rect 4344 24948 4396 24954
rect 4344 24890 4396 24896
rect 4816 24818 4844 25706
rect 5552 25498 5580 25842
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 3988 23322 4016 23666
rect 4172 23526 4200 24210
rect 4816 23730 4844 24754
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4908 24138 4936 24550
rect 5552 24206 5580 25434
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5644 24206 5672 24754
rect 5736 24342 5764 26386
rect 5816 26376 5868 26382
rect 5816 26318 5868 26324
rect 5724 24336 5776 24342
rect 5724 24278 5776 24284
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 4896 24132 4948 24138
rect 4896 24074 4948 24080
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4160 23520 4212 23526
rect 4160 23462 4212 23468
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 4528 23180 4580 23186
rect 4528 23122 4580 23128
rect 3884 23112 3936 23118
rect 3884 23054 3936 23060
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3896 19990 3924 23054
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 3988 21010 4016 21626
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 4264 19446 4292 20742
rect 4252 19440 4304 19446
rect 4252 19382 4304 19388
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3516 17264 3568 17270
rect 3516 17206 3568 17212
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3436 16250 3464 16934
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3804 14385 3832 18158
rect 3896 16590 3924 19246
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3988 18329 4016 19110
rect 4264 18766 4292 19246
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 3974 18320 4030 18329
rect 3974 18255 4030 18264
rect 4068 18284 4120 18290
rect 3988 18222 4016 18255
rect 4068 18226 4120 18232
rect 3976 18216 4028 18222
rect 4080 18193 4108 18226
rect 3976 18158 4028 18164
rect 4066 18184 4122 18193
rect 4066 18119 4122 18128
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 4080 16114 4108 18119
rect 4264 17814 4292 18702
rect 4356 18426 4384 21422
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4540 18306 4568 23122
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4632 22098 4660 22986
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4724 22234 4752 22578
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4620 22092 4672 22098
rect 4620 22034 4672 22040
rect 4816 20602 4844 23666
rect 4908 23089 4936 24074
rect 5736 24018 5764 24278
rect 5644 23990 5764 24018
rect 5644 23526 5672 23990
rect 5828 23866 5856 26318
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 5814 23624 5870 23633
rect 5814 23559 5870 23568
rect 5828 23526 5856 23559
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 4894 23080 4950 23089
rect 4894 23015 4950 23024
rect 5540 22976 5592 22982
rect 5540 22918 5592 22924
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 5000 20942 5028 22374
rect 5448 21616 5500 21622
rect 5448 21558 5500 21564
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 4804 20596 4856 20602
rect 4804 20538 4856 20544
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4712 18352 4764 18358
rect 4540 18278 4660 18306
rect 4712 18294 4764 18300
rect 4252 17808 4304 17814
rect 4252 17750 4304 17756
rect 4632 16289 4660 18278
rect 4724 16454 4752 18294
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4816 17270 4844 17614
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4618 16280 4674 16289
rect 4618 16215 4674 16224
rect 4908 16153 4936 18566
rect 5092 18426 5120 21286
rect 5460 21078 5488 21558
rect 5448 21072 5500 21078
rect 5448 21014 5500 21020
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 16590 5212 17682
rect 5368 17338 5396 19382
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5460 17134 5488 19178
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 4894 16144 4950 16153
rect 4068 16108 4120 16114
rect 5276 16114 5304 17002
rect 5460 16674 5488 17070
rect 5368 16646 5488 16674
rect 5368 16522 5396 16646
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 4894 16079 4950 16088
rect 5264 16108 5316 16114
rect 4068 16050 4120 16056
rect 5264 16050 5316 16056
rect 5276 15026 5304 16050
rect 5368 16046 5396 16458
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5368 15162 5396 15982
rect 5460 15502 5488 16526
rect 5552 16522 5580 22918
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5828 21554 5856 22374
rect 5920 21622 5948 26454
rect 6656 26450 6684 27950
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 6644 26444 6696 26450
rect 6644 26386 6696 26392
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6092 25152 6144 25158
rect 6092 25094 6144 25100
rect 6104 24886 6132 25094
rect 6092 24880 6144 24886
rect 6092 24822 6144 24828
rect 6104 23798 6132 24822
rect 6552 24676 6604 24682
rect 6552 24618 6604 24624
rect 6092 23792 6144 23798
rect 6092 23734 6144 23740
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 6012 22438 6040 23598
rect 6368 23588 6420 23594
rect 6368 23530 6420 23536
rect 6380 22642 6408 23530
rect 6564 23186 6592 24618
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6656 22778 6684 23666
rect 6840 23050 6868 25638
rect 7024 25158 7052 27338
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7012 25152 7064 25158
rect 7012 25094 7064 25100
rect 7300 24886 7328 25638
rect 7288 24880 7340 24886
rect 7288 24822 7340 24828
rect 7392 24614 7420 25774
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 6828 23044 6880 23050
rect 6828 22986 6880 22992
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6644 22568 6696 22574
rect 6748 22556 6776 22714
rect 6696 22528 6776 22556
rect 6644 22510 6696 22516
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 6184 21956 6236 21962
rect 6184 21898 6236 21904
rect 6196 21690 6224 21898
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6748 21622 6776 21830
rect 5908 21616 5960 21622
rect 5908 21558 5960 21564
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6748 21146 6776 21422
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6552 21004 6604 21010
rect 6552 20946 6604 20952
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5644 18290 5672 19654
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5736 18170 5764 19926
rect 6276 19780 6328 19786
rect 6276 19722 6328 19728
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 5920 18290 5948 18702
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5644 18142 5764 18170
rect 5644 17678 5672 18142
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5644 15638 5672 17614
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 5632 15632 5684 15638
rect 5632 15574 5684 15580
rect 5448 15496 5500 15502
rect 5736 15473 5764 17546
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5448 15438 5500 15444
rect 5722 15464 5778 15473
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5276 14618 5304 14962
rect 5460 14929 5488 15438
rect 5722 15399 5778 15408
rect 5446 14920 5502 14929
rect 5446 14855 5502 14864
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 3790 14376 3846 14385
rect 3790 14311 3846 14320
rect 5828 12345 5856 15914
rect 5920 14482 5948 17138
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6104 15502 6132 16730
rect 6196 15570 6224 19450
rect 6288 18426 6316 19722
rect 6380 19718 6408 20402
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6380 19378 6408 19654
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6288 16658 6316 18158
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6472 17542 6500 18022
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6564 17202 6592 20946
rect 6932 19310 6960 22714
rect 7012 22704 7064 22710
rect 7392 22681 7420 24550
rect 7012 22646 7064 22652
rect 7378 22672 7434 22681
rect 7024 21146 7052 22646
rect 7378 22607 7434 22616
rect 7104 22568 7156 22574
rect 7156 22528 7236 22556
rect 7104 22510 7156 22516
rect 7208 22094 7236 22528
rect 7208 22066 7328 22094
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7024 20466 7052 21082
rect 7116 20602 7144 21558
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7116 18698 7144 19314
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6288 16561 6316 16594
rect 6274 16552 6330 16561
rect 6274 16487 6330 16496
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 6012 13530 6040 15302
rect 6380 15026 6408 16458
rect 6458 16008 6514 16017
rect 6458 15943 6460 15952
rect 6512 15943 6514 15952
rect 6460 15914 6512 15920
rect 6564 15586 6592 16594
rect 6472 15558 6592 15586
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6472 13297 6500 15558
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6564 14890 6592 15438
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6656 14618 6684 18634
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6840 17490 6868 17546
rect 6840 17462 6960 17490
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6748 16182 6776 17070
rect 6736 16176 6788 16182
rect 6736 16118 6788 16124
rect 6748 15978 6776 16118
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6748 13938 6776 15438
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6840 14074 6868 15098
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6932 13462 6960 17462
rect 7024 17338 7052 18362
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7208 16590 7236 21286
rect 7300 20330 7328 22066
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7392 20602 7420 22034
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 7484 18714 7512 27406
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7668 24342 7696 26862
rect 7760 26382 7788 26930
rect 7748 26376 7800 26382
rect 7748 26318 7800 26324
rect 7852 26042 7880 28698
rect 7944 28558 7972 32438
rect 8036 31890 8064 33254
rect 8174 33212 8482 33221
rect 8174 33210 8180 33212
rect 8236 33210 8260 33212
rect 8316 33210 8340 33212
rect 8396 33210 8420 33212
rect 8476 33210 8482 33212
rect 8236 33158 8238 33210
rect 8418 33158 8420 33210
rect 8174 33156 8180 33158
rect 8236 33156 8260 33158
rect 8316 33156 8340 33158
rect 8396 33156 8420 33158
rect 8476 33156 8482 33158
rect 8174 33147 8482 33156
rect 9416 32774 9444 33458
rect 9404 32768 9456 32774
rect 9404 32710 9456 32716
rect 15398 32668 15706 32677
rect 15398 32666 15404 32668
rect 15460 32666 15484 32668
rect 15540 32666 15564 32668
rect 15620 32666 15644 32668
rect 15700 32666 15706 32668
rect 15460 32614 15462 32666
rect 15642 32614 15644 32666
rect 15398 32612 15404 32614
rect 15460 32612 15484 32614
rect 15540 32612 15564 32614
rect 15620 32612 15644 32614
rect 15700 32612 15706 32614
rect 15398 32603 15706 32612
rect 9036 32360 9088 32366
rect 9036 32302 9088 32308
rect 8174 32124 8482 32133
rect 8174 32122 8180 32124
rect 8236 32122 8260 32124
rect 8316 32122 8340 32124
rect 8396 32122 8420 32124
rect 8476 32122 8482 32124
rect 8236 32070 8238 32122
rect 8418 32070 8420 32122
rect 8174 32068 8180 32070
rect 8236 32068 8260 32070
rect 8316 32068 8340 32070
rect 8396 32068 8420 32070
rect 8476 32068 8482 32070
rect 8174 32059 8482 32068
rect 8024 31884 8076 31890
rect 8024 31826 8076 31832
rect 8036 31278 8064 31826
rect 8024 31272 8076 31278
rect 8024 31214 8076 31220
rect 8036 30734 8064 31214
rect 8174 31036 8482 31045
rect 8174 31034 8180 31036
rect 8236 31034 8260 31036
rect 8316 31034 8340 31036
rect 8396 31034 8420 31036
rect 8476 31034 8482 31036
rect 8236 30982 8238 31034
rect 8418 30982 8420 31034
rect 8174 30980 8180 30982
rect 8236 30980 8260 30982
rect 8316 30980 8340 30982
rect 8396 30980 8420 30982
rect 8476 30980 8482 30982
rect 8174 30971 8482 30980
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 8036 30054 8064 30670
rect 8024 30048 8076 30054
rect 8024 29990 8076 29996
rect 8036 29510 8064 29990
rect 8174 29948 8482 29957
rect 8174 29946 8180 29948
rect 8236 29946 8260 29948
rect 8316 29946 8340 29948
rect 8396 29946 8420 29948
rect 8476 29946 8482 29948
rect 8236 29894 8238 29946
rect 8418 29894 8420 29946
rect 8174 29892 8180 29894
rect 8236 29892 8260 29894
rect 8316 29892 8340 29894
rect 8396 29892 8420 29894
rect 8476 29892 8482 29894
rect 8174 29883 8482 29892
rect 8024 29504 8076 29510
rect 8024 29446 8076 29452
rect 8036 29102 8064 29446
rect 8024 29096 8076 29102
rect 8024 29038 8076 29044
rect 8760 29028 8812 29034
rect 8760 28970 8812 28976
rect 8174 28860 8482 28869
rect 8174 28858 8180 28860
rect 8236 28858 8260 28860
rect 8316 28858 8340 28860
rect 8396 28858 8420 28860
rect 8476 28858 8482 28860
rect 8236 28806 8238 28858
rect 8418 28806 8420 28858
rect 8174 28804 8180 28806
rect 8236 28804 8260 28806
rect 8316 28804 8340 28806
rect 8396 28804 8420 28806
rect 8476 28804 8482 28806
rect 8174 28795 8482 28804
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 7944 28150 7972 28494
rect 8024 28416 8076 28422
rect 8024 28358 8076 28364
rect 7932 28144 7984 28150
rect 7932 28086 7984 28092
rect 7944 27334 7972 28086
rect 7932 27328 7984 27334
rect 7932 27270 7984 27276
rect 7944 26450 7972 27270
rect 8036 26994 8064 28358
rect 8772 27946 8800 28970
rect 8852 28416 8904 28422
rect 8852 28358 8904 28364
rect 8760 27940 8812 27946
rect 8760 27882 8812 27888
rect 8174 27772 8482 27781
rect 8174 27770 8180 27772
rect 8236 27770 8260 27772
rect 8316 27770 8340 27772
rect 8396 27770 8420 27772
rect 8476 27770 8482 27772
rect 8236 27718 8238 27770
rect 8418 27718 8420 27770
rect 8174 27716 8180 27718
rect 8236 27716 8260 27718
rect 8316 27716 8340 27718
rect 8396 27716 8420 27718
rect 8476 27716 8482 27718
rect 8174 27707 8482 27716
rect 8576 27464 8628 27470
rect 8576 27406 8628 27412
rect 8024 26988 8076 26994
rect 8024 26930 8076 26936
rect 8588 26790 8616 27406
rect 8576 26784 8628 26790
rect 8576 26726 8628 26732
rect 8174 26684 8482 26693
rect 8174 26682 8180 26684
rect 8236 26682 8260 26684
rect 8316 26682 8340 26684
rect 8396 26682 8420 26684
rect 8476 26682 8482 26684
rect 8236 26630 8238 26682
rect 8418 26630 8420 26682
rect 8174 26628 8180 26630
rect 8236 26628 8260 26630
rect 8316 26628 8340 26630
rect 8396 26628 8420 26630
rect 8476 26628 8482 26630
rect 8174 26619 8482 26628
rect 8024 26512 8076 26518
rect 8024 26454 8076 26460
rect 7932 26444 7984 26450
rect 7932 26386 7984 26392
rect 8036 26234 8064 26454
rect 7944 26206 8064 26234
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7944 25362 7972 26206
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8174 25596 8482 25605
rect 8174 25594 8180 25596
rect 8236 25594 8260 25596
rect 8316 25594 8340 25596
rect 8396 25594 8420 25596
rect 8476 25594 8482 25596
rect 8236 25542 8238 25594
rect 8418 25542 8420 25594
rect 8174 25540 8180 25542
rect 8236 25540 8260 25542
rect 8316 25540 8340 25542
rect 8396 25540 8420 25542
rect 8476 25540 8482 25542
rect 8174 25531 8482 25540
rect 7932 25356 7984 25362
rect 7932 25298 7984 25304
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 7656 24336 7708 24342
rect 7656 24278 7708 24284
rect 7852 24206 7880 25230
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 8036 24290 8064 25162
rect 8174 24508 8482 24517
rect 8174 24506 8180 24508
rect 8236 24506 8260 24508
rect 8316 24506 8340 24508
rect 8396 24506 8420 24508
rect 8476 24506 8482 24508
rect 8236 24454 8238 24506
rect 8418 24454 8420 24506
rect 8174 24452 8180 24454
rect 8236 24452 8260 24454
rect 8316 24452 8340 24454
rect 8396 24452 8420 24454
rect 8476 24452 8482 24454
rect 8174 24443 8482 24452
rect 8114 24304 8170 24313
rect 8036 24262 8114 24290
rect 8114 24239 8116 24248
rect 8168 24239 8170 24248
rect 8116 24210 8168 24216
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7576 23322 7604 24142
rect 8588 23662 8616 25842
rect 8668 25696 8720 25702
rect 8668 25638 8720 25644
rect 8680 24818 8708 25638
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8772 24342 8800 24686
rect 8760 24336 8812 24342
rect 8760 24278 8812 24284
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7564 23044 7616 23050
rect 7616 23004 7696 23032
rect 7564 22986 7616 22992
rect 7668 22710 7696 23004
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7656 22704 7708 22710
rect 7656 22646 7708 22652
rect 7668 21962 7696 22646
rect 7760 22574 7788 22714
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7656 21956 7708 21962
rect 7656 21898 7708 21904
rect 7668 21078 7696 21898
rect 7656 21072 7708 21078
rect 7656 21014 7708 21020
rect 7668 20466 7696 21014
rect 7852 20534 7880 23530
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 22778 8064 23462
rect 8174 23420 8482 23429
rect 8174 23418 8180 23420
rect 8236 23418 8260 23420
rect 8316 23418 8340 23420
rect 8396 23418 8420 23420
rect 8476 23418 8482 23420
rect 8236 23366 8238 23418
rect 8418 23366 8420 23418
rect 8174 23364 8180 23366
rect 8236 23364 8260 23366
rect 8316 23364 8340 23366
rect 8396 23364 8420 23366
rect 8476 23364 8482 23366
rect 8174 23355 8482 23364
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 8174 22332 8482 22341
rect 8174 22330 8180 22332
rect 8236 22330 8260 22332
rect 8316 22330 8340 22332
rect 8396 22330 8420 22332
rect 8476 22330 8482 22332
rect 8236 22278 8238 22330
rect 8418 22278 8420 22330
rect 8174 22276 8180 22278
rect 8236 22276 8260 22278
rect 8316 22276 8340 22278
rect 8396 22276 8420 22278
rect 8476 22276 8482 22278
rect 8174 22267 8482 22276
rect 8024 21956 8076 21962
rect 7944 21916 8024 21944
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7944 20058 7972 21916
rect 8024 21898 8076 21904
rect 8174 21244 8482 21253
rect 8174 21242 8180 21244
rect 8236 21242 8260 21244
rect 8316 21242 8340 21244
rect 8396 21242 8420 21244
rect 8476 21242 8482 21244
rect 8236 21190 8238 21242
rect 8418 21190 8420 21242
rect 8174 21188 8180 21190
rect 8236 21188 8260 21190
rect 8316 21188 8340 21190
rect 8396 21188 8420 21190
rect 8476 21188 8482 21190
rect 8174 21179 8482 21188
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8174 20156 8482 20165
rect 8174 20154 8180 20156
rect 8236 20154 8260 20156
rect 8316 20154 8340 20156
rect 8396 20154 8420 20156
rect 8476 20154 8482 20156
rect 8236 20102 8238 20154
rect 8418 20102 8420 20154
rect 8174 20100 8180 20102
rect 8236 20100 8260 20102
rect 8316 20100 8340 20102
rect 8396 20100 8420 20102
rect 8476 20100 8482 20102
rect 8174 20091 8482 20100
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7668 19446 7696 19722
rect 7656 19440 7708 19446
rect 7656 19382 7708 19388
rect 8174 19068 8482 19077
rect 8174 19066 8180 19068
rect 8236 19066 8260 19068
rect 8316 19066 8340 19068
rect 8396 19066 8420 19068
rect 8476 19066 8482 19068
rect 8236 19014 8238 19066
rect 8418 19014 8420 19066
rect 8174 19012 8180 19014
rect 8236 19012 8260 19014
rect 8316 19012 8340 19014
rect 8396 19012 8420 19014
rect 8476 19012 8482 19014
rect 8174 19003 8482 19012
rect 7392 18686 7512 18714
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 18358 7328 18566
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 7392 17066 7420 18686
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7208 16114 7236 16526
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7484 15026 7512 18566
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8174 17980 8482 17989
rect 8174 17978 8180 17980
rect 8236 17978 8260 17980
rect 8316 17978 8340 17980
rect 8396 17978 8420 17980
rect 8476 17978 8482 17980
rect 8236 17926 8238 17978
rect 8418 17926 8420 17978
rect 8174 17924 8180 17926
rect 8236 17924 8260 17926
rect 8316 17924 8340 17926
rect 8396 17924 8420 17926
rect 8476 17924 8482 17926
rect 8174 17915 8482 17924
rect 8588 17338 8616 18022
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8174 16892 8482 16901
rect 8174 16890 8180 16892
rect 8236 16890 8260 16892
rect 8316 16890 8340 16892
rect 8396 16890 8420 16892
rect 8476 16890 8482 16892
rect 8236 16838 8238 16890
rect 8418 16838 8420 16890
rect 8174 16836 8180 16838
rect 8236 16836 8260 16838
rect 8316 16836 8340 16838
rect 8396 16836 8420 16838
rect 8476 16836 8482 16838
rect 8174 16827 8482 16836
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6458 13288 6514 13297
rect 6458 13223 6514 13232
rect 7484 12850 7512 14962
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 5814 12336 5870 12345
rect 5814 12271 5870 12280
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1596 10305 1624 10610
rect 1582 10296 1638 10305
rect 1582 10231 1584 10240
rect 1636 10231 1638 10240
rect 1584 10202 1636 10208
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3252 9178 3280 9318
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4865 1532 4966
rect 1490 4856 1546 4865
rect 1490 4791 1546 4800
rect 1688 2446 1716 8774
rect 7576 7478 7604 15302
rect 7944 15026 7972 15846
rect 8174 15804 8482 15813
rect 8174 15802 8180 15804
rect 8236 15802 8260 15804
rect 8316 15802 8340 15804
rect 8396 15802 8420 15804
rect 8476 15802 8482 15804
rect 8236 15750 8238 15802
rect 8418 15750 8420 15802
rect 8174 15748 8180 15750
rect 8236 15748 8260 15750
rect 8316 15748 8340 15750
rect 8396 15748 8420 15750
rect 8476 15748 8482 15750
rect 8174 15739 8482 15748
rect 8298 15600 8354 15609
rect 8298 15535 8300 15544
rect 8352 15535 8354 15544
rect 8300 15506 8352 15512
rect 8680 15434 8708 17478
rect 8772 17134 8800 20198
rect 8864 18578 8892 28358
rect 9048 27985 9076 32302
rect 15398 31580 15706 31589
rect 15398 31578 15404 31580
rect 15460 31578 15484 31580
rect 15540 31578 15564 31580
rect 15620 31578 15644 31580
rect 15700 31578 15706 31580
rect 15460 31526 15462 31578
rect 15642 31526 15644 31578
rect 15398 31524 15404 31526
rect 15460 31524 15484 31526
rect 15540 31524 15564 31526
rect 15620 31524 15644 31526
rect 15700 31524 15706 31526
rect 15398 31515 15706 31524
rect 15398 30492 15706 30501
rect 15398 30490 15404 30492
rect 15460 30490 15484 30492
rect 15540 30490 15564 30492
rect 15620 30490 15644 30492
rect 15700 30490 15706 30492
rect 15460 30438 15462 30490
rect 15642 30438 15644 30490
rect 15398 30436 15404 30438
rect 15460 30436 15484 30438
rect 15540 30436 15564 30438
rect 15620 30436 15644 30438
rect 15700 30436 15706 30438
rect 15398 30427 15706 30436
rect 14372 30252 14424 30258
rect 14372 30194 14424 30200
rect 14384 29646 14412 30194
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 14568 29714 14596 30126
rect 15200 30048 15252 30054
rect 15200 29990 15252 29996
rect 15212 29850 15240 29990
rect 15200 29844 15252 29850
rect 15200 29786 15252 29792
rect 14556 29708 14608 29714
rect 14556 29650 14608 29656
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 9588 29504 9640 29510
rect 9588 29446 9640 29452
rect 9600 28422 9628 29446
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9588 28416 9640 28422
rect 9588 28358 9640 28364
rect 9128 28144 9180 28150
rect 9128 28086 9180 28092
rect 9034 27976 9090 27985
rect 9034 27911 9090 27920
rect 8944 27328 8996 27334
rect 8944 27270 8996 27276
rect 8956 27130 8984 27270
rect 8944 27124 8996 27130
rect 8944 27066 8996 27072
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 8956 26382 8984 26862
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 8944 25288 8996 25294
rect 8944 25230 8996 25236
rect 8956 21894 8984 25230
rect 9048 23866 9076 27911
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 9140 23746 9168 28086
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 9416 26382 9444 27406
rect 9600 27334 9628 28358
rect 9692 27946 9720 28562
rect 14384 28558 14412 29582
rect 14568 28626 14596 29650
rect 16488 29572 16540 29578
rect 16488 29514 16540 29520
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 15398 29404 15706 29413
rect 15398 29402 15404 29404
rect 15460 29402 15484 29404
rect 15540 29402 15564 29404
rect 15620 29402 15644 29404
rect 15700 29402 15706 29404
rect 15460 29350 15462 29402
rect 15642 29350 15644 29402
rect 15398 29348 15404 29350
rect 15460 29348 15484 29350
rect 15540 29348 15564 29350
rect 15620 29348 15644 29350
rect 15700 29348 15706 29350
rect 15398 29339 15706 29348
rect 14556 28620 14608 28626
rect 14556 28562 14608 28568
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 9680 27940 9732 27946
rect 9680 27882 9732 27888
rect 9692 27538 9720 27882
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 14384 27470 14412 28494
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15304 27538 15332 28358
rect 15398 28316 15706 28325
rect 15398 28314 15404 28316
rect 15460 28314 15484 28316
rect 15540 28314 15564 28316
rect 15620 28314 15644 28316
rect 15700 28314 15706 28316
rect 15460 28262 15462 28314
rect 15642 28262 15644 28314
rect 15398 28260 15404 28262
rect 15460 28260 15484 28262
rect 15540 28260 15564 28262
rect 15620 28260 15644 28262
rect 15700 28260 15706 28262
rect 15398 28251 15706 28260
rect 15292 27532 15344 27538
rect 15292 27474 15344 27480
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 15764 27334 15792 29446
rect 16500 29306 16528 29514
rect 16488 29300 16540 29306
rect 16488 29242 16540 29248
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16776 27674 16804 27814
rect 16764 27668 16816 27674
rect 16764 27610 16816 27616
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 10876 27328 10928 27334
rect 10876 27270 10928 27276
rect 15752 27328 15804 27334
rect 15752 27270 15804 27276
rect 9956 27056 10008 27062
rect 9956 26998 10008 27004
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9232 25906 9260 26250
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9416 25498 9444 26318
rect 9876 26314 9904 26794
rect 9968 26450 9996 26998
rect 10888 26586 10916 27270
rect 15398 27228 15706 27237
rect 15398 27226 15404 27228
rect 15460 27226 15484 27228
rect 15540 27226 15564 27228
rect 15620 27226 15644 27228
rect 15700 27226 15706 27228
rect 15460 27174 15462 27226
rect 15642 27174 15644 27226
rect 15398 27172 15404 27174
rect 15460 27172 15484 27174
rect 15540 27172 15564 27174
rect 15620 27172 15644 27174
rect 15700 27172 15706 27174
rect 15398 27163 15706 27172
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 15292 26988 15344 26994
rect 15292 26930 15344 26936
rect 13820 26852 13872 26858
rect 13820 26794 13872 26800
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 12256 26512 12308 26518
rect 12256 26454 12308 26460
rect 9956 26444 10008 26450
rect 9956 26386 10008 26392
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 9220 25424 9272 25430
rect 9220 25366 9272 25372
rect 9232 24750 9260 25366
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9692 24698 9720 24822
rect 9692 24670 9812 24698
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9692 24206 9720 24550
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9048 23718 9168 23746
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8864 18550 8984 18578
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 8772 15570 8800 16526
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 12782 7788 14214
rect 7852 13802 7880 14758
rect 7944 14482 7972 14962
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 8036 14006 8064 14758
rect 8174 14716 8482 14725
rect 8174 14714 8180 14716
rect 8236 14714 8260 14716
rect 8316 14714 8340 14716
rect 8396 14714 8420 14716
rect 8476 14714 8482 14716
rect 8236 14662 8238 14714
rect 8418 14662 8420 14714
rect 8174 14660 8180 14662
rect 8236 14660 8260 14662
rect 8316 14660 8340 14662
rect 8396 14660 8420 14662
rect 8476 14660 8482 14662
rect 8174 14651 8482 14660
rect 8300 14544 8352 14550
rect 8298 14512 8300 14521
rect 8352 14512 8354 14521
rect 8298 14447 8354 14456
rect 8680 14414 8708 15370
rect 8864 14618 8892 15846
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8956 14550 8984 18550
rect 9048 16726 9076 23718
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9140 20602 9168 23598
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9140 19242 9168 19858
rect 9128 19236 9180 19242
rect 9128 19178 9180 19184
rect 9140 17202 9168 19178
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 9232 16590 9260 18022
rect 9324 17785 9352 23802
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9692 23118 9720 23462
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9784 22710 9812 24670
rect 9876 23322 9904 26250
rect 9968 25974 9996 26386
rect 11060 26376 11112 26382
rect 11060 26318 11112 26324
rect 11072 26042 11100 26318
rect 11060 26036 11112 26042
rect 11060 25978 11112 25984
rect 9956 25968 10008 25974
rect 9956 25910 10008 25916
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 10888 25498 10916 25774
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 10980 25294 11008 25842
rect 12268 25838 12296 26454
rect 12544 26314 12572 26726
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 12256 25832 12308 25838
rect 12256 25774 12308 25780
rect 11072 25362 11100 25774
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 9968 24410 9996 25230
rect 10980 24818 11008 25230
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 10704 24274 10732 24550
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10968 24132 11020 24138
rect 10968 24074 11020 24080
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 9416 20942 9444 21558
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9692 19514 9720 21898
rect 9784 20534 9812 22646
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9876 19854 9904 23258
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 10152 21962 10180 22918
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9310 17776 9366 17785
rect 9310 17711 9366 17720
rect 9600 17678 9628 19110
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9784 17610 9812 19654
rect 10244 19378 10272 19790
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9126 16280 9182 16289
rect 9126 16215 9182 16224
rect 9140 15706 9168 16215
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9232 15586 9260 16526
rect 9140 15558 9260 15586
rect 9508 15570 9536 16594
rect 9876 16250 9904 18634
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10244 18426 10272 18566
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10336 17202 10364 20946
rect 10428 20058 10456 21490
rect 10980 21418 11008 24074
rect 11164 23338 11192 25366
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 11164 23310 11284 23338
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11072 22710 11100 23054
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 11164 22506 11192 23122
rect 11152 22500 11204 22506
rect 11152 22442 11204 22448
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10796 20466 10824 20742
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10796 19854 10824 20402
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10796 16658 10824 17138
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9496 15564 9548 15570
rect 9140 15502 9168 15558
rect 9496 15506 9548 15512
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8758 13968 8814 13977
rect 7932 13932 7984 13938
rect 8758 13903 8760 13912
rect 7932 13874 7984 13880
rect 8812 13903 8814 13912
rect 8760 13874 8812 13880
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7944 13326 7972 13874
rect 9232 13870 9260 15438
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14414 9720 14758
rect 9876 14482 9904 16186
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9968 14618 9996 16118
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 8036 13394 8064 13806
rect 8174 13628 8482 13637
rect 8174 13626 8180 13628
rect 8236 13626 8260 13628
rect 8316 13626 8340 13628
rect 8396 13626 8420 13628
rect 8476 13626 8482 13628
rect 8236 13574 8238 13626
rect 8418 13574 8420 13626
rect 8174 13572 8180 13574
rect 8236 13572 8260 13574
rect 8316 13572 8340 13574
rect 8396 13572 8420 13574
rect 8476 13572 8482 13574
rect 8174 13563 8482 13572
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 8036 13190 8064 13330
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 9692 12986 9720 14350
rect 10060 12986 10088 16390
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10612 15706 10640 15982
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 14006 10456 15438
rect 10704 14958 10732 15982
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10612 14618 10640 14894
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10600 14272 10652 14278
rect 10704 14226 10732 14894
rect 10652 14220 10732 14226
rect 10600 14214 10732 14220
rect 10612 14198 10732 14214
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 10428 13530 10456 13942
rect 10704 13870 10732 14198
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7944 6798 7972 12582
rect 8174 12540 8482 12549
rect 8174 12538 8180 12540
rect 8236 12538 8260 12540
rect 8316 12538 8340 12540
rect 8396 12538 8420 12540
rect 8476 12538 8482 12540
rect 8236 12486 8238 12538
rect 8418 12486 8420 12538
rect 8174 12484 8180 12486
rect 8236 12484 8260 12486
rect 8316 12484 8340 12486
rect 8396 12484 8420 12486
rect 8476 12484 8482 12486
rect 8174 12475 8482 12484
rect 10796 12442 10824 16594
rect 10888 15502 10916 19314
rect 11072 17882 11100 19722
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10888 14550 10916 15098
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10980 12918 11008 15642
rect 11072 15638 11100 17070
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 11164 12850 11192 21830
rect 11256 19922 11284 23310
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11348 19514 11376 22170
rect 11440 20466 11468 25094
rect 11704 24404 11756 24410
rect 11704 24346 11756 24352
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 11624 19718 11652 21830
rect 11716 21554 11744 24346
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11808 21690 11836 23054
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11796 21548 11848 21554
rect 11796 21490 11848 21496
rect 11808 20602 11836 21490
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11796 20392 11848 20398
rect 11796 20334 11848 20340
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 18902 11376 19110
rect 11336 18896 11388 18902
rect 11336 18838 11388 18844
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11256 16658 11284 18362
rect 11348 18222 11376 18566
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11348 16454 11376 18158
rect 11440 17882 11468 19382
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11532 18630 11560 18838
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11532 17814 11560 18566
rect 11716 18290 11744 19314
rect 11808 18970 11836 20334
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11900 18766 11928 19314
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11624 17270 11652 18022
rect 11716 17678 11744 18226
rect 11980 18148 12032 18154
rect 11980 18090 12032 18096
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11808 14074 11836 17546
rect 11900 17542 11928 17750
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11992 16046 12020 18090
rect 12084 17105 12112 25638
rect 12164 25424 12216 25430
rect 12164 25366 12216 25372
rect 12268 25378 12296 25774
rect 12544 25770 12572 26250
rect 12532 25764 12584 25770
rect 12532 25706 12584 25712
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 12622 25392 12678 25401
rect 12176 23050 12204 25366
rect 12268 25362 12388 25378
rect 12268 25356 12400 25362
rect 12268 25350 12348 25356
rect 12268 24818 12296 25350
rect 12622 25327 12624 25336
rect 12348 25298 12400 25304
rect 12676 25327 12678 25336
rect 12624 25298 12676 25304
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12636 24886 12664 25162
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 12624 24880 12676 24886
rect 12624 24822 12676 24828
rect 12912 24818 12940 25094
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12268 24206 12296 24754
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12164 23044 12216 23050
rect 12164 22986 12216 22992
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 21962 12480 22374
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12544 21010 12572 22578
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12360 19922 12756 19938
rect 12360 19916 12768 19922
rect 12360 19910 12716 19916
rect 12360 19446 12388 19910
rect 12716 19858 12768 19864
rect 12532 19780 12584 19786
rect 12532 19722 12584 19728
rect 12544 19514 12572 19722
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12912 19310 12940 24754
rect 13280 24274 13308 25434
rect 13372 24410 13400 26318
rect 13452 26308 13504 26314
rect 13452 26250 13504 26256
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 13176 23792 13228 23798
rect 13176 23734 13228 23740
rect 13084 23656 13136 23662
rect 13084 23598 13136 23604
rect 12992 21344 13044 21350
rect 13096 21332 13124 23598
rect 13188 23118 13216 23734
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13188 22642 13216 23054
rect 13280 22778 13308 24210
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13188 21690 13216 22578
rect 13372 22098 13400 24210
rect 13464 23730 13492 26250
rect 13832 25906 13860 26794
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 14200 25974 14228 26726
rect 14476 26382 14504 26930
rect 14556 26920 14608 26926
rect 14556 26862 14608 26868
rect 14464 26376 14516 26382
rect 14464 26318 14516 26324
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 14476 25838 14504 26318
rect 14464 25832 14516 25838
rect 14464 25774 14516 25780
rect 13636 25764 13688 25770
rect 13636 25706 13688 25712
rect 13544 25696 13596 25702
rect 13544 25638 13596 25644
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 13360 22092 13412 22098
rect 13464 22094 13492 23530
rect 13556 22794 13584 25638
rect 13648 24177 13676 25706
rect 13728 24676 13780 24682
rect 13728 24618 13780 24624
rect 13634 24168 13690 24177
rect 13634 24103 13690 24112
rect 13648 23186 13676 24103
rect 13740 23594 13768 24618
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13728 23588 13780 23594
rect 13728 23530 13780 23536
rect 13636 23180 13688 23186
rect 13636 23122 13688 23128
rect 13556 22766 13676 22794
rect 13464 22066 13584 22094
rect 13360 22034 13412 22040
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13044 21304 13124 21332
rect 12992 21286 13044 21292
rect 13004 19378 13032 21286
rect 13556 20942 13584 22066
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 13188 19174 13216 20198
rect 13556 19718 13584 20266
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13096 17542 13124 18294
rect 13188 18290 13216 19110
rect 13280 18766 13308 19246
rect 13372 18834 13400 19654
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13280 18358 13308 18702
rect 13372 18630 13400 18770
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12070 17096 12126 17105
rect 12070 17031 12126 17040
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12268 16182 12296 17002
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16182 12756 16934
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11440 13802 11468 14010
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 8174 11452 8482 11461
rect 8174 11450 8180 11452
rect 8236 11450 8260 11452
rect 8316 11450 8340 11452
rect 8396 11450 8420 11452
rect 8476 11450 8482 11452
rect 8236 11398 8238 11450
rect 8418 11398 8420 11450
rect 8174 11396 8180 11398
rect 8236 11396 8260 11398
rect 8316 11396 8340 11398
rect 8396 11396 8420 11398
rect 8476 11396 8482 11398
rect 8174 11387 8482 11396
rect 11900 11150 11928 12786
rect 11992 11830 12020 15982
rect 13004 15570 13032 15982
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12084 12850 12112 15438
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12544 14958 12572 15030
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12268 11898 12296 14758
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12360 14074 12388 14214
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12348 13932 12400 13938
rect 12452 13920 12480 14282
rect 12400 13892 12480 13920
rect 12348 13874 12400 13880
rect 12452 13530 12480 13892
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12622 12880 12678 12889
rect 12622 12815 12624 12824
rect 12676 12815 12678 12824
rect 12624 12786 12676 12792
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 12636 11762 12664 12174
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12820 11354 12848 14350
rect 13096 12170 13124 17478
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 13280 11898 13308 16662
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13372 14414 13400 15438
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13556 12850 13584 13738
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13464 12434 13492 12718
rect 13372 12406 13492 12434
rect 13372 12306 13400 12406
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13372 11354 13400 12242
rect 13556 12238 13584 12786
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11801 13584 12038
rect 13542 11792 13598 11801
rect 13542 11727 13598 11736
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 8174 10364 8482 10373
rect 8174 10362 8180 10364
rect 8236 10362 8260 10364
rect 8316 10362 8340 10364
rect 8396 10362 8420 10364
rect 8476 10362 8482 10364
rect 8236 10310 8238 10362
rect 8418 10310 8420 10362
rect 8174 10308 8180 10310
rect 8236 10308 8260 10310
rect 8316 10308 8340 10310
rect 8396 10308 8420 10310
rect 8476 10308 8482 10310
rect 8174 10299 8482 10308
rect 8174 9276 8482 9285
rect 8174 9274 8180 9276
rect 8236 9274 8260 9276
rect 8316 9274 8340 9276
rect 8396 9274 8420 9276
rect 8476 9274 8482 9276
rect 8236 9222 8238 9274
rect 8418 9222 8420 9274
rect 8174 9220 8180 9222
rect 8236 9220 8260 9222
rect 8316 9220 8340 9222
rect 8396 9220 8420 9222
rect 8476 9220 8482 9222
rect 8174 9211 8482 9220
rect 8174 8188 8482 8197
rect 8174 8186 8180 8188
rect 8236 8186 8260 8188
rect 8316 8186 8340 8188
rect 8396 8186 8420 8188
rect 8476 8186 8482 8188
rect 8236 8134 8238 8186
rect 8418 8134 8420 8186
rect 8174 8132 8180 8134
rect 8236 8132 8260 8134
rect 8316 8132 8340 8134
rect 8396 8132 8420 8134
rect 8476 8132 8482 8134
rect 8174 8123 8482 8132
rect 8174 7100 8482 7109
rect 8174 7098 8180 7100
rect 8236 7098 8260 7100
rect 8316 7098 8340 7100
rect 8396 7098 8420 7100
rect 8476 7098 8482 7100
rect 8236 7046 8238 7098
rect 8418 7046 8420 7098
rect 8174 7044 8180 7046
rect 8236 7044 8260 7046
rect 8316 7044 8340 7046
rect 8396 7044 8420 7046
rect 8476 7044 8482 7046
rect 8174 7035 8482 7044
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 8174 6012 8482 6021
rect 8174 6010 8180 6012
rect 8236 6010 8260 6012
rect 8316 6010 8340 6012
rect 8396 6010 8420 6012
rect 8476 6010 8482 6012
rect 8236 5958 8238 6010
rect 8418 5958 8420 6010
rect 8174 5956 8180 5958
rect 8236 5956 8260 5958
rect 8316 5956 8340 5958
rect 8396 5956 8420 5958
rect 8476 5956 8482 5958
rect 8174 5947 8482 5956
rect 8174 4924 8482 4933
rect 8174 4922 8180 4924
rect 8236 4922 8260 4924
rect 8316 4922 8340 4924
rect 8396 4922 8420 4924
rect 8476 4922 8482 4924
rect 8236 4870 8238 4922
rect 8418 4870 8420 4922
rect 8174 4868 8180 4870
rect 8236 4868 8260 4870
rect 8316 4868 8340 4870
rect 8396 4868 8420 4870
rect 8476 4868 8482 4870
rect 8174 4859 8482 4868
rect 13648 4146 13676 22766
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13740 21962 13768 22714
rect 13728 21956 13780 21962
rect 13728 21898 13780 21904
rect 13924 20058 13952 23666
rect 14108 22710 14136 24550
rect 14476 24410 14504 25774
rect 14568 25430 14596 26862
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 15108 26444 15160 26450
rect 15108 26386 15160 26392
rect 14556 25424 14608 25430
rect 14556 25366 14608 25372
rect 14660 25294 14688 26386
rect 15016 26308 15068 26314
rect 15016 26250 15068 26256
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14936 24410 14964 24686
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14660 23798 14688 24142
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 15028 23050 15056 26250
rect 15016 23044 15068 23050
rect 14936 23004 15016 23032
rect 14936 22778 14964 23004
rect 15016 22986 15068 22992
rect 15120 22794 15148 26386
rect 15304 25922 15332 26930
rect 15764 26382 15792 26998
rect 15936 26920 15988 26926
rect 15936 26862 15988 26868
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15844 26376 15896 26382
rect 15844 26318 15896 26324
rect 15398 26140 15706 26149
rect 15398 26138 15404 26140
rect 15460 26138 15484 26140
rect 15540 26138 15564 26140
rect 15620 26138 15644 26140
rect 15700 26138 15706 26140
rect 15460 26086 15462 26138
rect 15642 26086 15644 26138
rect 15398 26084 15404 26086
rect 15460 26084 15484 26086
rect 15540 26084 15564 26086
rect 15620 26084 15644 26086
rect 15700 26084 15706 26086
rect 15398 26075 15706 26084
rect 15856 26042 15884 26318
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15384 25968 15436 25974
rect 15304 25916 15384 25922
rect 15948 25922 15976 26862
rect 17236 26586 17264 33458
rect 19444 33114 19472 33458
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 27344 33312 27396 33318
rect 27344 33254 27396 33260
rect 22622 33212 22930 33221
rect 22622 33210 22628 33212
rect 22684 33210 22708 33212
rect 22764 33210 22788 33212
rect 22844 33210 22868 33212
rect 22924 33210 22930 33212
rect 22684 33158 22686 33210
rect 22866 33158 22868 33210
rect 22622 33156 22628 33158
rect 22684 33156 22708 33158
rect 22764 33156 22788 33158
rect 22844 33156 22868 33158
rect 22924 33156 22930 33158
rect 22622 33147 22930 33156
rect 19432 33108 19484 33114
rect 19432 33050 19484 33056
rect 18696 32904 18748 32910
rect 18696 32846 18748 32852
rect 18708 31754 18736 32846
rect 24308 32768 24360 32774
rect 24308 32710 24360 32716
rect 22622 32124 22930 32133
rect 22622 32122 22628 32124
rect 22684 32122 22708 32124
rect 22764 32122 22788 32124
rect 22844 32122 22868 32124
rect 22924 32122 22930 32124
rect 22684 32070 22686 32122
rect 22866 32070 22868 32122
rect 22622 32068 22628 32070
rect 22684 32068 22708 32070
rect 22764 32068 22788 32070
rect 22844 32068 22868 32070
rect 22924 32068 22930 32070
rect 22622 32059 22930 32068
rect 18616 31726 18736 31754
rect 18616 29578 18644 31726
rect 22622 31036 22930 31045
rect 22622 31034 22628 31036
rect 22684 31034 22708 31036
rect 22764 31034 22788 31036
rect 22844 31034 22868 31036
rect 22924 31034 22930 31036
rect 22684 30982 22686 31034
rect 22866 30982 22868 31034
rect 22622 30980 22628 30982
rect 22684 30980 22708 30982
rect 22764 30980 22788 30982
rect 22844 30980 22868 30982
rect 22924 30980 22930 30982
rect 22622 30971 22930 30980
rect 19524 30252 19576 30258
rect 19524 30194 19576 30200
rect 19536 29714 19564 30194
rect 20720 30048 20772 30054
rect 20720 29990 20772 29996
rect 20732 29714 20760 29990
rect 22622 29948 22930 29957
rect 22622 29946 22628 29948
rect 22684 29946 22708 29948
rect 22764 29946 22788 29948
rect 22844 29946 22868 29948
rect 22924 29946 22930 29948
rect 22684 29894 22686 29946
rect 22866 29894 22868 29946
rect 22622 29892 22628 29894
rect 22684 29892 22708 29894
rect 22764 29892 22788 29894
rect 22844 29892 22868 29894
rect 22924 29892 22930 29894
rect 22622 29883 22930 29892
rect 19524 29708 19576 29714
rect 19524 29650 19576 29656
rect 20720 29708 20772 29714
rect 20720 29650 20772 29656
rect 18604 29572 18656 29578
rect 18604 29514 18656 29520
rect 18052 28960 18104 28966
rect 18052 28902 18104 28908
rect 17776 28552 17828 28558
rect 17776 28494 17828 28500
rect 17788 28014 17816 28494
rect 18064 28422 18092 28902
rect 18616 28762 18644 29514
rect 19248 29504 19300 29510
rect 19248 29446 19300 29452
rect 19260 29170 19288 29446
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19536 29102 19564 29650
rect 24124 29640 24176 29646
rect 24124 29582 24176 29588
rect 20628 29572 20680 29578
rect 20628 29514 20680 29520
rect 19524 29096 19576 29102
rect 19524 29038 19576 29044
rect 18604 28756 18656 28762
rect 18604 28698 18656 28704
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 18064 28218 18092 28358
rect 18052 28212 18104 28218
rect 18052 28154 18104 28160
rect 17776 28008 17828 28014
rect 17776 27950 17828 27956
rect 17788 27674 17816 27950
rect 18064 27826 18092 28154
rect 18616 28150 18644 28698
rect 20352 28416 20404 28422
rect 20352 28358 20404 28364
rect 20364 28150 20392 28358
rect 20640 28218 20668 29514
rect 24136 29306 24164 29582
rect 24124 29300 24176 29306
rect 24124 29242 24176 29248
rect 21732 29096 21784 29102
rect 21732 29038 21784 29044
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 20352 28144 20404 28150
rect 20352 28086 20404 28092
rect 19340 27940 19392 27946
rect 19340 27882 19392 27888
rect 18064 27798 18184 27826
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 18052 27396 18104 27402
rect 18052 27338 18104 27344
rect 18064 27130 18092 27338
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 17684 27056 17736 27062
rect 17684 26998 17736 27004
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 17224 26580 17276 26586
rect 17224 26522 17276 26528
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 15304 25910 15436 25916
rect 15304 25894 15424 25910
rect 15856 25894 15976 25922
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 15212 24750 15240 25230
rect 15398 25052 15706 25061
rect 15398 25050 15404 25052
rect 15460 25050 15484 25052
rect 15540 25050 15564 25052
rect 15620 25050 15644 25052
rect 15700 25050 15706 25052
rect 15460 24998 15462 25050
rect 15642 24998 15644 25050
rect 15398 24996 15404 24998
rect 15460 24996 15484 24998
rect 15540 24996 15564 24998
rect 15620 24996 15644 24998
rect 15700 24996 15706 24998
rect 15398 24987 15706 24996
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15856 24614 15884 25894
rect 17052 25838 17080 26182
rect 17040 25832 17092 25838
rect 17040 25774 17092 25780
rect 16672 25764 16724 25770
rect 16672 25706 16724 25712
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15200 24132 15252 24138
rect 15200 24074 15252 24080
rect 15212 23866 15240 24074
rect 15200 23860 15252 23866
rect 15200 23802 15252 23808
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 15028 22766 15148 22794
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14016 19514 14044 20402
rect 14108 19854 14136 21830
rect 14476 20602 14504 22374
rect 14936 22094 14964 22714
rect 15028 22522 15056 22766
rect 15028 22494 15148 22522
rect 14936 22066 15056 22094
rect 15028 21962 15056 22066
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 15028 21554 15056 21898
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14384 19514 14412 19654
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13740 13190 13768 18634
rect 14568 18630 14596 19654
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14568 18193 14596 18566
rect 14660 18426 14688 20810
rect 14740 19712 14792 19718
rect 15120 19666 15148 22494
rect 15212 20942 15240 23802
rect 15304 23304 15332 24142
rect 15398 23964 15706 23973
rect 15398 23962 15404 23964
rect 15460 23962 15484 23964
rect 15540 23962 15564 23964
rect 15620 23962 15644 23964
rect 15700 23962 15706 23964
rect 15460 23910 15462 23962
rect 15642 23910 15644 23962
rect 15398 23908 15404 23910
rect 15460 23908 15484 23910
rect 15540 23908 15564 23910
rect 15620 23908 15644 23910
rect 15700 23908 15706 23910
rect 15398 23899 15706 23908
rect 15384 23316 15436 23322
rect 15304 23276 15384 23304
rect 15384 23258 15436 23264
rect 15398 22876 15706 22885
rect 15398 22874 15404 22876
rect 15460 22874 15484 22876
rect 15540 22874 15564 22876
rect 15620 22874 15644 22876
rect 15700 22874 15706 22876
rect 15460 22822 15462 22874
rect 15642 22822 15644 22874
rect 15398 22820 15404 22822
rect 15460 22820 15484 22822
rect 15540 22820 15564 22822
rect 15620 22820 15644 22822
rect 15700 22820 15706 22822
rect 15398 22811 15706 22820
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15304 21486 15332 22510
rect 15856 22094 15884 24550
rect 15948 23186 15976 25094
rect 16040 24954 16068 25230
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 16040 22642 16068 24890
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16132 23662 16160 24550
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16212 23044 16264 23050
rect 16212 22986 16264 22992
rect 16028 22636 16080 22642
rect 16080 22596 16160 22624
rect 16028 22578 16080 22584
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 16040 22098 16068 22374
rect 15856 22066 15976 22094
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15398 21788 15706 21797
rect 15398 21786 15404 21788
rect 15460 21786 15484 21788
rect 15540 21786 15564 21788
rect 15620 21786 15644 21788
rect 15700 21786 15706 21788
rect 15460 21734 15462 21786
rect 15642 21734 15644 21786
rect 15398 21732 15404 21734
rect 15460 21732 15484 21734
rect 15540 21732 15564 21734
rect 15620 21732 15644 21734
rect 15700 21732 15706 21734
rect 15398 21723 15706 21732
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15764 21350 15792 21490
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20602 15240 20742
rect 15398 20700 15706 20709
rect 15398 20698 15404 20700
rect 15460 20698 15484 20700
rect 15540 20698 15564 20700
rect 15620 20698 15644 20700
rect 15700 20698 15706 20700
rect 15460 20646 15462 20698
rect 15642 20646 15644 20698
rect 15398 20644 15404 20646
rect 15460 20644 15484 20646
rect 15540 20644 15564 20646
rect 15620 20644 15644 20646
rect 15700 20644 15706 20646
rect 15398 20635 15706 20644
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15580 19990 15608 20198
rect 15856 20097 15884 21898
rect 15842 20088 15898 20097
rect 15842 20023 15898 20032
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 14740 19654 14792 19660
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14752 18290 14780 19654
rect 14936 19638 15148 19666
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14554 18184 14610 18193
rect 14554 18119 14610 18128
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14108 16697 14136 18022
rect 14094 16688 14150 16697
rect 14094 16623 14150 16632
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 16250 14320 16390
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13832 14346 13860 15302
rect 13924 14618 13952 15370
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 14016 13938 14044 14758
rect 14384 14550 14412 16050
rect 14752 15978 14780 18226
rect 14936 17241 14964 19638
rect 15398 19612 15706 19621
rect 15398 19610 15404 19612
rect 15460 19610 15484 19612
rect 15540 19610 15564 19612
rect 15620 19610 15644 19612
rect 15700 19610 15706 19612
rect 15460 19558 15462 19610
rect 15642 19558 15644 19610
rect 15398 19556 15404 19558
rect 15460 19556 15484 19558
rect 15540 19556 15564 19558
rect 15620 19556 15644 19558
rect 15700 19556 15706 19558
rect 15398 19547 15706 19556
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 14922 17232 14978 17241
rect 14922 17167 14978 17176
rect 15028 16658 15056 19314
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15120 17649 15148 18770
rect 15398 18524 15706 18533
rect 15398 18522 15404 18524
rect 15460 18522 15484 18524
rect 15540 18522 15564 18524
rect 15620 18522 15644 18524
rect 15700 18522 15706 18524
rect 15460 18470 15462 18522
rect 15642 18470 15644 18522
rect 15398 18468 15404 18470
rect 15460 18468 15484 18470
rect 15540 18468 15564 18470
rect 15620 18468 15644 18470
rect 15700 18468 15706 18470
rect 15398 18459 15706 18468
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15200 17672 15252 17678
rect 15106 17640 15162 17649
rect 15200 17614 15252 17620
rect 15106 17575 15162 17584
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13924 13258 13952 13806
rect 14384 13326 14412 14214
rect 14752 13870 14780 14554
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 13740 12782 13768 13126
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 14292 12646 14320 13126
rect 14384 12918 14412 13262
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14752 12442 14780 13806
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14844 11898 14872 16594
rect 15212 16454 15240 17614
rect 15304 17270 15332 17818
rect 15948 17746 15976 22066
rect 16028 22092 16080 22098
rect 16028 22034 16080 22040
rect 16132 21146 16160 22596
rect 16224 22234 16252 22986
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16316 22642 16344 22918
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16580 22568 16632 22574
rect 16684 22556 16712 25706
rect 17052 24750 17080 25774
rect 17408 25288 17460 25294
rect 17406 25256 17408 25265
rect 17460 25256 17462 25265
rect 17406 25191 17462 25200
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17040 24744 17092 24750
rect 17040 24686 17092 24692
rect 17052 24206 17080 24686
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 17328 23662 17356 24754
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 17224 23248 17276 23254
rect 17224 23190 17276 23196
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16632 22528 16712 22556
rect 16580 22510 16632 22516
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16592 22094 16620 22374
rect 16684 22166 16712 22528
rect 16672 22160 16724 22166
rect 16672 22102 16724 22108
rect 16408 22066 16620 22094
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16316 21622 16344 21966
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 16408 21554 16436 22066
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16408 20466 16436 21490
rect 16500 20942 16528 21966
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16500 20806 16528 20878
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16500 20466 16528 20742
rect 16776 20618 16804 22918
rect 17052 22778 17080 23190
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17236 22681 17264 23190
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 17222 22672 17278 22681
rect 17222 22607 17278 22616
rect 17132 22500 17184 22506
rect 17132 22442 17184 22448
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17052 21010 17080 22034
rect 17144 21622 17172 22442
rect 17328 22094 17356 22714
rect 17420 22642 17448 23054
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17408 22094 17460 22098
rect 17328 22092 17460 22094
rect 17328 22066 17408 22092
rect 17408 22034 17460 22040
rect 17132 21616 17184 21622
rect 17132 21558 17184 21564
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 16592 20590 16804 20618
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 16488 20460 16540 20466
rect 16488 20402 16540 20408
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16500 19689 16528 19858
rect 16592 19825 16620 20590
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 16776 20262 16804 20470
rect 17052 20398 17080 20946
rect 17040 20392 17092 20398
rect 17040 20334 17092 20340
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16578 19816 16634 19825
rect 16578 19751 16634 19760
rect 16486 19680 16542 19689
rect 16486 19615 16542 19624
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16040 18465 16068 18702
rect 16026 18456 16082 18465
rect 16026 18391 16082 18400
rect 16488 18420 16540 18426
rect 16040 18154 16068 18391
rect 16488 18362 16540 18368
rect 16028 18148 16080 18154
rect 16028 18090 16080 18096
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15398 17436 15706 17445
rect 15398 17434 15404 17436
rect 15460 17434 15484 17436
rect 15540 17434 15564 17436
rect 15620 17434 15644 17436
rect 15700 17434 15706 17436
rect 15460 17382 15462 17434
rect 15642 17382 15644 17434
rect 15398 17380 15404 17382
rect 15460 17380 15484 17382
rect 15540 17380 15564 17382
rect 15620 17380 15644 17382
rect 15700 17380 15706 17382
rect 15398 17371 15706 17380
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 15212 15502 15240 16390
rect 15398 16348 15706 16357
rect 15398 16346 15404 16348
rect 15460 16346 15484 16348
rect 15540 16346 15564 16348
rect 15620 16346 15644 16348
rect 15700 16346 15706 16348
rect 15460 16294 15462 16346
rect 15642 16294 15644 16346
rect 15398 16292 15404 16294
rect 15460 16292 15484 16294
rect 15540 16292 15564 16294
rect 15620 16292 15644 16294
rect 15700 16292 15706 16294
rect 15398 16283 15706 16292
rect 15764 16182 15792 16390
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 16132 15910 16160 16390
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15212 15162 15240 15438
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15304 15094 15332 15846
rect 15398 15260 15706 15269
rect 15398 15258 15404 15260
rect 15460 15258 15484 15260
rect 15540 15258 15564 15260
rect 15620 15258 15644 15260
rect 15700 15258 15706 15260
rect 15460 15206 15462 15258
rect 15642 15206 15644 15258
rect 15398 15204 15404 15206
rect 15460 15204 15484 15206
rect 15540 15204 15564 15206
rect 15620 15204 15644 15206
rect 15700 15204 15706 15206
rect 15398 15195 15706 15204
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15304 13394 15332 15030
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15398 14172 15706 14181
rect 15398 14170 15404 14172
rect 15460 14170 15484 14172
rect 15540 14170 15564 14172
rect 15620 14170 15644 14172
rect 15700 14170 15706 14172
rect 15460 14118 15462 14170
rect 15642 14118 15644 14170
rect 15398 14116 15404 14118
rect 15460 14116 15484 14118
rect 15540 14116 15564 14118
rect 15620 14116 15644 14118
rect 15700 14116 15706 14118
rect 15398 14107 15706 14116
rect 15764 13394 15792 14418
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16040 14074 16068 14350
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15398 13084 15706 13093
rect 15398 13082 15404 13084
rect 15460 13082 15484 13084
rect 15540 13082 15564 13084
rect 15620 13082 15644 13084
rect 15700 13082 15706 13084
rect 15460 13030 15462 13082
rect 15642 13030 15644 13082
rect 15398 13028 15404 13030
rect 15460 13028 15484 13030
rect 15540 13028 15564 13030
rect 15620 13028 15644 13030
rect 15700 13028 15706 13030
rect 15398 13019 15706 13028
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 15028 12434 15056 12650
rect 15856 12434 15884 13670
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15028 12406 15148 12434
rect 15856 12406 15976 12434
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 15120 11558 15148 12406
rect 15398 11996 15706 12005
rect 15398 11994 15404 11996
rect 15460 11994 15484 11996
rect 15540 11994 15564 11996
rect 15620 11994 15644 11996
rect 15700 11994 15706 11996
rect 15460 11942 15462 11994
rect 15642 11942 15644 11994
rect 15398 11940 15404 11942
rect 15460 11940 15484 11942
rect 15540 11940 15564 11942
rect 15620 11940 15644 11942
rect 15700 11940 15706 11942
rect 15398 11931 15706 11940
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 11150 15148 11494
rect 15948 11234 15976 12406
rect 16040 11370 16068 13262
rect 16224 11830 16252 17818
rect 16500 17202 16528 18362
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16500 16726 16528 17138
rect 16592 17134 16620 19751
rect 16776 19242 16804 20198
rect 17052 19310 17080 20334
rect 17144 19854 17172 21014
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17420 19786 17448 21286
rect 17408 19780 17460 19786
rect 17408 19722 17460 19728
rect 17420 19514 17448 19722
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17328 18698 17356 19110
rect 17316 18692 17368 18698
rect 17316 18634 17368 18640
rect 17512 17218 17540 26930
rect 17696 26586 17724 26998
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17684 26580 17736 26586
rect 17684 26522 17736 26528
rect 17696 26382 17724 26522
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17592 25356 17644 25362
rect 17592 25298 17644 25304
rect 17604 24750 17632 25298
rect 17592 24744 17644 24750
rect 17592 24686 17644 24692
rect 17604 24410 17632 24686
rect 17592 24404 17644 24410
rect 17592 24346 17644 24352
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 17338 17632 17478
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17512 17190 17632 17218
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16592 16794 16620 17070
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16592 16538 16620 16594
rect 17222 16552 17278 16561
rect 16592 16510 16804 16538
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 16046 16344 16390
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16500 14414 16528 15642
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16578 14376 16634 14385
rect 16578 14311 16634 14320
rect 16592 13938 16620 14311
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16394 12200 16450 12209
rect 16394 12135 16396 12144
rect 16448 12135 16450 12144
rect 16396 12106 16448 12112
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16040 11342 16252 11370
rect 15948 11218 16068 11234
rect 15948 11212 16080 11218
rect 15948 11206 16028 11212
rect 16028 11154 16080 11160
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15398 10908 15706 10917
rect 15398 10906 15404 10908
rect 15460 10906 15484 10908
rect 15540 10906 15564 10908
rect 15620 10906 15644 10908
rect 15700 10906 15706 10908
rect 15460 10854 15462 10906
rect 15642 10854 15644 10906
rect 15398 10852 15404 10854
rect 15460 10852 15484 10854
rect 15540 10852 15564 10854
rect 15620 10852 15644 10854
rect 15700 10852 15706 10854
rect 15398 10843 15706 10852
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 9926 13860 10406
rect 15764 9926 15792 11086
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 16040 10810 16068 11018
rect 16224 11014 16252 11342
rect 16592 11234 16620 13194
rect 16684 11354 16712 15370
rect 16776 15026 16804 16510
rect 17222 16487 17278 16496
rect 17236 16046 17264 16487
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16776 12442 16804 14962
rect 17500 14952 17552 14958
rect 17498 14920 17500 14929
rect 17552 14920 17554 14929
rect 17498 14855 17554 14864
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 14074 17172 14350
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17328 14074 17356 14282
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17052 13258 17080 13466
rect 17314 13288 17370 13297
rect 17040 13252 17092 13258
rect 17314 13223 17370 13232
rect 17040 13194 17092 13200
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16868 11694 16896 12378
rect 16960 12102 16988 12922
rect 17328 12918 17356 13223
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 17052 11762 17080 12718
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17144 12170 17172 12582
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 17604 11898 17632 17190
rect 17696 12434 17724 26318
rect 17880 25838 17908 26726
rect 18156 26518 18184 27798
rect 19352 27554 19380 27882
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19352 27526 19472 27554
rect 19628 27538 19656 27814
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 18144 26512 18196 26518
rect 18144 26454 18196 26460
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17776 25764 17828 25770
rect 17776 25706 17828 25712
rect 17788 25294 17816 25706
rect 17776 25288 17828 25294
rect 17776 25230 17828 25236
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17788 21418 17816 22578
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17880 20534 17908 25774
rect 18052 25424 18104 25430
rect 18052 25366 18104 25372
rect 18064 23322 18092 25366
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18156 24138 18184 24550
rect 18144 24132 18196 24138
rect 18144 24074 18196 24080
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18050 23080 18106 23089
rect 17960 23044 18012 23050
rect 18050 23015 18052 23024
rect 17960 22986 18012 22992
rect 18104 23015 18106 23024
rect 18052 22986 18104 22992
rect 17972 21690 18000 22986
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17788 18714 17816 20198
rect 17880 20058 17908 20470
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17788 18686 17908 18714
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17788 18057 17816 18566
rect 17774 18048 17830 18057
rect 17774 17983 17830 17992
rect 17880 16794 17908 18686
rect 17972 17270 18000 19314
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17960 17128 18012 17134
rect 18064 17082 18092 18634
rect 18012 17076 18092 17082
rect 17960 17070 18092 17076
rect 17972 17054 18092 17070
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17788 16674 17816 16730
rect 17788 16646 17908 16674
rect 17880 16590 17908 16646
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17972 13172 18000 13942
rect 18156 13841 18184 24074
rect 18248 19530 18276 27406
rect 19444 27402 19472 27526
rect 19616 27532 19668 27538
rect 19616 27474 19668 27480
rect 19432 27396 19484 27402
rect 19432 27338 19484 27344
rect 20720 26852 20772 26858
rect 20720 26794 20772 26800
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 18972 26512 19024 26518
rect 18972 26454 19024 26460
rect 18328 25832 18380 25838
rect 18328 25774 18380 25780
rect 18340 25498 18368 25774
rect 18328 25492 18380 25498
rect 18328 25434 18380 25440
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18340 25265 18368 25298
rect 18326 25256 18382 25265
rect 18326 25191 18382 25200
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18340 24206 18368 24754
rect 18512 24676 18564 24682
rect 18512 24618 18564 24624
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18340 23730 18368 24142
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18340 21978 18368 23258
rect 18418 23216 18474 23225
rect 18418 23151 18474 23160
rect 18432 22545 18460 23151
rect 18418 22536 18474 22545
rect 18418 22471 18420 22480
rect 18472 22471 18474 22480
rect 18420 22442 18472 22448
rect 18432 22411 18460 22442
rect 18524 22438 18552 24618
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18420 22094 18472 22098
rect 18524 22094 18552 22374
rect 18616 22098 18644 23258
rect 18420 22092 18552 22094
rect 18472 22066 18552 22092
rect 18604 22092 18656 22098
rect 18420 22034 18472 22040
rect 18604 22034 18656 22040
rect 18340 21950 18552 21978
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18340 20398 18368 21422
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18340 19990 18368 20334
rect 18328 19984 18380 19990
rect 18432 19961 18460 20742
rect 18328 19926 18380 19932
rect 18418 19952 18474 19961
rect 18418 19887 18474 19896
rect 18248 19502 18368 19530
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 18248 18766 18276 19382
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18248 16998 18276 18702
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18248 16658 18276 16934
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18142 13832 18198 13841
rect 18142 13767 18198 13776
rect 17972 13144 18092 13172
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17696 12406 17816 12434
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 17408 11688 17460 11694
rect 17408 11630 17460 11636
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16592 11206 16712 11234
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16224 10674 16252 10950
rect 16592 10742 16620 11018
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16224 10266 16252 10610
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16684 10198 16712 11206
rect 17420 11014 17448 11630
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17052 10538 17080 10950
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17040 10532 17092 10538
rect 17040 10474 17092 10480
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 8174 3836 8482 3845
rect 8174 3834 8180 3836
rect 8236 3834 8260 3836
rect 8316 3834 8340 3836
rect 8396 3834 8420 3836
rect 8476 3834 8482 3836
rect 8236 3782 8238 3834
rect 8418 3782 8420 3834
rect 8174 3780 8180 3782
rect 8236 3780 8260 3782
rect 8316 3780 8340 3782
rect 8396 3780 8420 3782
rect 8476 3780 8482 3782
rect 8174 3771 8482 3780
rect 8174 2748 8482 2757
rect 8174 2746 8180 2748
rect 8236 2746 8260 2748
rect 8316 2746 8340 2748
rect 8396 2746 8420 2748
rect 8476 2746 8482 2748
rect 8236 2694 8238 2746
rect 8418 2694 8420 2746
rect 8174 2692 8180 2694
rect 8236 2692 8260 2694
rect 8316 2692 8340 2694
rect 8396 2692 8420 2694
rect 8476 2692 8482 2694
rect 8174 2683 8482 2692
rect 13832 2582 13860 9862
rect 15398 9820 15706 9829
rect 15398 9818 15404 9820
rect 15460 9818 15484 9820
rect 15540 9818 15564 9820
rect 15620 9818 15644 9820
rect 15700 9818 15706 9820
rect 15460 9766 15462 9818
rect 15642 9766 15644 9818
rect 15398 9764 15404 9766
rect 15460 9764 15484 9766
rect 15540 9764 15564 9766
rect 15620 9764 15644 9766
rect 15700 9764 15706 9766
rect 15398 9755 15706 9764
rect 17604 9722 17632 10678
rect 17696 10606 17724 11562
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 8838 16344 9318
rect 17604 8906 17632 9658
rect 17788 9450 17816 12406
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 11150 17908 11698
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17880 10742 17908 10950
rect 17972 10810 18000 12922
rect 18064 11354 18092 13144
rect 18340 12986 18368 19502
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18432 18358 18460 18702
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18420 17604 18472 17610
rect 18420 17546 18472 17552
rect 18432 16590 18460 17546
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18524 14482 18552 21950
rect 18708 21554 18736 25094
rect 18788 24812 18840 24818
rect 18840 24772 18920 24800
rect 18788 24754 18840 24760
rect 18892 23186 18920 24772
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18892 21865 18920 23122
rect 18984 23118 19012 26454
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19628 25906 19656 26318
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 19800 25696 19852 25702
rect 19800 25638 19852 25644
rect 19616 25356 19668 25362
rect 19616 25298 19668 25304
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18878 21856 18934 21865
rect 18878 21791 18934 21800
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18708 20942 18736 21490
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18616 17814 18644 18770
rect 18694 18456 18750 18465
rect 18694 18391 18750 18400
rect 18708 18358 18736 18391
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18708 17814 18736 18158
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18604 16516 18656 16522
rect 18604 16458 18656 16464
rect 18616 15706 18644 16458
rect 18696 16040 18748 16046
rect 18694 16008 18696 16017
rect 18748 16008 18750 16017
rect 18694 15943 18750 15952
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18800 15570 18828 19450
rect 18892 19378 18920 21791
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 19076 18290 19104 24210
rect 19168 23526 19196 24754
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 19168 21962 19196 23462
rect 19536 23322 19564 25162
rect 19628 24750 19656 25298
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19628 24274 19656 24686
rect 19616 24268 19668 24274
rect 19616 24210 19668 24216
rect 19628 23662 19656 24210
rect 19720 23746 19748 25230
rect 19812 24886 19840 25638
rect 20088 25226 20116 26726
rect 20352 26444 20404 26450
rect 20352 26386 20404 26392
rect 20364 25838 20392 26386
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20456 26042 20484 26318
rect 20628 26240 20680 26246
rect 20628 26182 20680 26188
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20444 25900 20496 25906
rect 20444 25842 20496 25848
rect 20352 25832 20404 25838
rect 20352 25774 20404 25780
rect 20364 25294 20392 25774
rect 20456 25294 20484 25842
rect 20352 25288 20404 25294
rect 20352 25230 20404 25236
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 19800 24880 19852 24886
rect 19800 24822 19852 24828
rect 19892 24608 19944 24614
rect 19892 24550 19944 24556
rect 19904 23769 19932 24550
rect 19890 23760 19946 23769
rect 19720 23718 19840 23746
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 19156 21956 19208 21962
rect 19156 21898 19208 21904
rect 19260 21486 19288 22986
rect 19340 22024 19392 22030
rect 19338 21992 19340 22001
rect 19392 21992 19394 22001
rect 19338 21927 19394 21936
rect 19444 21729 19472 23190
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19430 21720 19486 21729
rect 19430 21655 19486 21664
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19168 20330 19196 21354
rect 19260 20618 19288 21422
rect 19444 21146 19472 21655
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19260 20602 19380 20618
rect 19260 20596 19392 20602
rect 19260 20590 19340 20596
rect 19340 20538 19392 20544
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19260 18737 19288 19654
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19246 18728 19302 18737
rect 19246 18663 19302 18672
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18984 16250 19012 18226
rect 19352 17610 19380 19382
rect 19444 19242 19472 19858
rect 19432 19236 19484 19242
rect 19432 19178 19484 19184
rect 19536 18426 19564 23122
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19628 21622 19656 21966
rect 19616 21616 19668 21622
rect 19616 21558 19668 21564
rect 19628 21078 19656 21558
rect 19616 21072 19668 21078
rect 19616 21014 19668 21020
rect 19616 19848 19668 19854
rect 19614 19816 19616 19825
rect 19668 19816 19670 19825
rect 19614 19751 19670 19760
rect 19720 19514 19748 22986
rect 19812 21486 19840 23718
rect 19890 23695 19946 23704
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19996 23118 20024 23598
rect 20088 23186 20116 25162
rect 20456 24070 20484 25230
rect 20640 24750 20668 26182
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20548 24313 20576 24550
rect 20534 24304 20590 24313
rect 20534 24239 20590 24248
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 20260 23588 20312 23594
rect 20260 23530 20312 23536
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20180 21690 20208 21830
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 20272 21010 20300 23530
rect 20732 23225 20760 26794
rect 20904 25832 20956 25838
rect 20904 25774 20956 25780
rect 20812 25764 20864 25770
rect 20812 25706 20864 25712
rect 20824 24721 20852 25706
rect 20810 24712 20866 24721
rect 20810 24647 20866 24656
rect 20718 23216 20774 23225
rect 20718 23151 20774 23160
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20352 22160 20404 22166
rect 20352 22102 20404 22108
rect 20364 21418 20392 22102
rect 20352 21412 20404 21418
rect 20352 21354 20404 21360
rect 20260 21004 20312 21010
rect 20260 20946 20312 20952
rect 20364 20942 20392 21354
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20456 20806 20484 23054
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20548 21146 20576 22918
rect 20732 22642 20760 23151
rect 20916 22778 20944 25774
rect 21548 25764 21600 25770
rect 21548 25706 21600 25712
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 21008 24070 21036 25298
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21468 25158 21496 25230
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 21456 25152 21508 25158
rect 21456 25094 21508 25100
rect 21284 24818 21312 25094
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21088 24744 21140 24750
rect 21088 24686 21140 24692
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 21100 23633 21128 24686
rect 21364 24200 21416 24206
rect 21362 24168 21364 24177
rect 21416 24168 21418 24177
rect 21362 24103 21418 24112
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21086 23624 21142 23633
rect 21086 23559 21142 23568
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20640 22234 20668 22374
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20640 22030 20668 22170
rect 20916 22166 20944 22714
rect 20904 22160 20956 22166
rect 20904 22102 20956 22108
rect 21008 22094 21036 23122
rect 21192 23118 21220 23666
rect 21468 23662 21496 25094
rect 21456 23656 21508 23662
rect 21456 23598 21508 23604
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21192 22438 21220 23054
rect 21364 23044 21416 23050
rect 21364 22986 21416 22992
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21284 22506 21312 22714
rect 21272 22500 21324 22506
rect 21272 22442 21324 22448
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 21088 22094 21140 22098
rect 21008 22092 21140 22094
rect 21008 22066 21088 22092
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 21008 21894 21036 22066
rect 21088 22034 21140 22040
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21100 21690 21128 21830
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 19890 19816 19946 19825
rect 19890 19751 19946 19760
rect 19904 19718 19932 19751
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19628 18902 19656 19246
rect 19616 18896 19668 18902
rect 19616 18838 19668 18844
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 18984 14521 19012 14894
rect 19260 14618 19288 15030
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19352 14550 19380 16662
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19444 15638 19472 15982
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19340 14544 19392 14550
rect 18970 14512 19026 14521
rect 18512 14476 18564 14482
rect 19340 14486 19392 14492
rect 18970 14447 19026 14456
rect 18512 14418 18564 14424
rect 19444 14396 19472 15098
rect 19536 14890 19564 15438
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19536 14414 19564 14826
rect 19352 14368 19472 14396
rect 19524 14408 19576 14414
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18524 14074 18552 14214
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18604 13252 18656 13258
rect 18604 13194 18656 13200
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 18616 12782 18644 13194
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 18156 10130 18184 12650
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18328 12368 18380 12374
rect 18328 12310 18380 12316
rect 18248 12102 18276 12310
rect 18340 12209 18368 12310
rect 18326 12200 18382 12209
rect 18326 12135 18382 12144
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18708 11898 18736 13942
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18616 9926 18644 10746
rect 18800 9926 18828 13126
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18984 12238 19012 12718
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 19352 10674 19380 14368
rect 19524 14350 19576 14356
rect 19628 14260 19656 18838
rect 19996 18834 20024 19314
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20272 17882 20300 18022
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20456 17678 20484 19858
rect 20628 19780 20680 19786
rect 20628 19722 20680 19728
rect 20640 17678 20668 19722
rect 20732 18766 20760 21422
rect 21100 21078 21128 21626
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21088 21072 21140 21078
rect 21088 21014 21140 21020
rect 21284 21010 21312 21286
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20916 20058 20944 20538
rect 21284 20398 21312 20946
rect 21376 20602 21404 22986
rect 21560 22094 21588 25706
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21652 23118 21680 24550
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21560 22066 21680 22094
rect 21652 21350 21680 22066
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21548 21072 21600 21078
rect 21546 21040 21548 21049
rect 21600 21040 21602 21049
rect 21546 20975 21602 20984
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20916 19854 20944 19994
rect 21284 19854 21312 20198
rect 20904 19848 20956 19854
rect 21272 19848 21324 19854
rect 20956 19808 21036 19836
rect 20904 19790 20956 19796
rect 21008 18970 21036 19808
rect 21272 19790 21324 19796
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21192 18766 21220 19110
rect 20720 18760 20772 18766
rect 21180 18760 21232 18766
rect 20720 18702 20772 18708
rect 21100 18720 21180 18748
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 19812 17338 19840 17614
rect 20456 17542 20484 17614
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 19800 17332 19852 17338
rect 19800 17274 19852 17280
rect 19706 16280 19762 16289
rect 19706 16215 19762 16224
rect 19720 16182 19748 16215
rect 19708 16176 19760 16182
rect 19708 16118 19760 16124
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20074 16008 20130 16017
rect 20074 15943 20130 15952
rect 20088 15570 20116 15943
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19444 14232 19656 14260
rect 19444 12442 19472 14232
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11665 19472 12038
rect 19536 11830 19564 12310
rect 19628 11898 19656 13670
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19524 11688 19576 11694
rect 19430 11656 19486 11665
rect 19524 11630 19576 11636
rect 19430 11591 19486 11600
rect 19536 11150 19564 11630
rect 19720 11218 19748 14894
rect 19812 14618 19840 15438
rect 20180 15162 20208 16118
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 14618 19932 14758
rect 19800 14612 19852 14618
rect 19800 14554 19852 14560
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 20272 14346 20300 15982
rect 20640 15706 20668 17614
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20732 15094 20760 17070
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20824 16266 20852 16594
rect 21008 16454 21036 17546
rect 21100 16658 21128 18720
rect 21180 18702 21232 18708
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21192 18426 21220 18566
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21192 18086 21220 18362
rect 21180 18080 21232 18086
rect 21232 18040 21312 18068
rect 21180 18022 21232 18028
rect 21178 17096 21234 17105
rect 21178 17031 21180 17040
rect 21232 17031 21234 17040
rect 21180 17002 21232 17008
rect 21192 16658 21220 17002
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 20824 16238 20944 16266
rect 20916 15609 20944 16238
rect 21100 15910 21128 16594
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 20902 15600 20958 15609
rect 20902 15535 20958 15544
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20824 14414 20852 14962
rect 20812 14408 20864 14414
rect 20864 14368 20944 14396
rect 20812 14350 20864 14356
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 20260 14340 20312 14346
rect 20260 14282 20312 14288
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19904 12850 19932 13262
rect 19996 12918 20024 13806
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 20180 11778 20208 14282
rect 20272 13938 20300 14282
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20272 12374 20300 13874
rect 20916 12434 20944 14368
rect 21008 14113 21036 15846
rect 21100 15162 21128 15846
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 21100 14464 21128 14962
rect 21180 14476 21232 14482
rect 21100 14436 21180 14464
rect 21180 14418 21232 14424
rect 20994 14104 21050 14113
rect 20994 14039 21050 14048
rect 21008 13938 21036 14039
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20916 12406 21036 12434
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20180 11762 20300 11778
rect 20180 11756 20312 11762
rect 20180 11750 20260 11756
rect 20260 11698 20312 11704
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19352 9994 19380 10610
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18418 9616 18474 9625
rect 18418 9551 18474 9560
rect 18432 9518 18460 9551
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 18708 9178 18736 9454
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 15398 8732 15706 8741
rect 15398 8730 15404 8732
rect 15460 8730 15484 8732
rect 15540 8730 15564 8732
rect 15620 8730 15644 8732
rect 15700 8730 15706 8732
rect 15460 8678 15462 8730
rect 15642 8678 15644 8730
rect 15398 8676 15404 8678
rect 15460 8676 15484 8678
rect 15540 8676 15564 8678
rect 15620 8676 15644 8678
rect 15700 8676 15706 8678
rect 15398 8667 15706 8676
rect 15398 7644 15706 7653
rect 15398 7642 15404 7644
rect 15460 7642 15484 7644
rect 15540 7642 15564 7644
rect 15620 7642 15644 7644
rect 15700 7642 15706 7644
rect 15460 7590 15462 7642
rect 15642 7590 15644 7642
rect 15398 7588 15404 7590
rect 15460 7588 15484 7590
rect 15540 7588 15564 7590
rect 15620 7588 15644 7590
rect 15700 7588 15706 7590
rect 15398 7579 15706 7588
rect 15398 6556 15706 6565
rect 15398 6554 15404 6556
rect 15460 6554 15484 6556
rect 15540 6554 15564 6556
rect 15620 6554 15644 6556
rect 15700 6554 15706 6556
rect 15460 6502 15462 6554
rect 15642 6502 15644 6554
rect 15398 6500 15404 6502
rect 15460 6500 15484 6502
rect 15540 6500 15564 6502
rect 15620 6500 15644 6502
rect 15700 6500 15706 6502
rect 15398 6491 15706 6500
rect 15398 5468 15706 5477
rect 15398 5466 15404 5468
rect 15460 5466 15484 5468
rect 15540 5466 15564 5468
rect 15620 5466 15644 5468
rect 15700 5466 15706 5468
rect 15460 5414 15462 5466
rect 15642 5414 15644 5466
rect 15398 5412 15404 5414
rect 15460 5412 15484 5414
rect 15540 5412 15564 5414
rect 15620 5412 15644 5414
rect 15700 5412 15706 5414
rect 15398 5403 15706 5412
rect 15398 4380 15706 4389
rect 15398 4378 15404 4380
rect 15460 4378 15484 4380
rect 15540 4378 15564 4380
rect 15620 4378 15644 4380
rect 15700 4378 15706 4380
rect 15460 4326 15462 4378
rect 15642 4326 15644 4378
rect 15398 4324 15404 4326
rect 15460 4324 15484 4326
rect 15540 4324 15564 4326
rect 15620 4324 15644 4326
rect 15700 4324 15706 4326
rect 15398 4315 15706 4324
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14292 3194 14320 4082
rect 15398 3292 15706 3301
rect 15398 3290 15404 3292
rect 15460 3290 15484 3292
rect 15540 3290 15564 3292
rect 15620 3290 15644 3292
rect 15700 3290 15706 3292
rect 15460 3238 15462 3290
rect 15642 3238 15644 3290
rect 15398 3236 15404 3238
rect 15460 3236 15484 3238
rect 15540 3236 15564 3238
rect 15620 3236 15644 3238
rect 15700 3236 15706 3238
rect 15398 3227 15706 3236
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 14292 2446 14320 3130
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 32 800 60 2246
rect 4540 800 4568 2382
rect 16316 2378 16344 8774
rect 17144 8634 17172 8842
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 18800 8498 18828 9862
rect 19904 9178 19932 11154
rect 20272 10062 20300 11698
rect 20364 10606 20392 12038
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 20444 10736 20496 10742
rect 20444 10678 20496 10684
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20272 9722 20300 9862
rect 20456 9722 20484 10678
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20732 9654 20760 11154
rect 21008 10470 21036 12406
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21100 11626 21128 12174
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 19892 9172 19944 9178
rect 19892 9114 19944 9120
rect 20272 9110 20300 9318
rect 21008 9178 21036 10406
rect 21100 10062 21128 11562
rect 21192 10810 21220 14418
rect 21284 14414 21312 18040
rect 21376 15162 21404 18634
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21638 15056 21694 15065
rect 21638 14991 21694 15000
rect 21652 14958 21680 14991
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21364 14272 21416 14278
rect 21416 14232 21496 14260
rect 21364 14214 21416 14220
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21376 11762 21404 12310
rect 21468 11762 21496 14232
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11286 21404 11494
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21192 10198 21220 10610
rect 21180 10192 21232 10198
rect 21180 10134 21232 10140
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20260 9104 20312 9110
rect 20260 9046 20312 9052
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19996 8634 20024 8842
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 19996 8362 20024 8570
rect 20272 8566 20300 9046
rect 21178 8936 21234 8945
rect 21178 8871 21234 8880
rect 21192 8838 21220 8871
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 20456 7886 20484 8774
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20548 7886 20576 8298
rect 21192 8294 21220 8774
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21192 8090 21220 8230
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20548 6866 20576 7822
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20916 7410 20944 7686
rect 21640 7472 21692 7478
rect 21640 7414 21692 7420
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 21652 7002 21680 7414
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19536 6458 19564 6734
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19720 5370 19748 6598
rect 21744 5370 21772 29038
rect 22622 28860 22930 28869
rect 22622 28858 22628 28860
rect 22684 28858 22708 28860
rect 22764 28858 22788 28860
rect 22844 28858 22868 28860
rect 22924 28858 22930 28860
rect 22684 28806 22686 28858
rect 22866 28806 22868 28858
rect 22622 28804 22628 28806
rect 22684 28804 22708 28806
rect 22764 28804 22788 28806
rect 22844 28804 22868 28806
rect 22924 28804 22930 28806
rect 22622 28795 22930 28804
rect 22622 27772 22930 27781
rect 22622 27770 22628 27772
rect 22684 27770 22708 27772
rect 22764 27770 22788 27772
rect 22844 27770 22868 27772
rect 22924 27770 22930 27772
rect 22684 27718 22686 27770
rect 22866 27718 22868 27770
rect 22622 27716 22628 27718
rect 22684 27716 22708 27718
rect 22764 27716 22788 27718
rect 22844 27716 22868 27718
rect 22924 27716 22930 27718
rect 22622 27707 22930 27716
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 23020 26852 23072 26858
rect 23020 26794 23072 26800
rect 22622 26684 22930 26693
rect 22622 26682 22628 26684
rect 22684 26682 22708 26684
rect 22764 26682 22788 26684
rect 22844 26682 22868 26684
rect 22924 26682 22930 26684
rect 22684 26630 22686 26682
rect 22866 26630 22868 26682
rect 22622 26628 22628 26630
rect 22684 26628 22708 26630
rect 22764 26628 22788 26630
rect 22844 26628 22868 26630
rect 22924 26628 22930 26630
rect 22622 26619 22930 26628
rect 22376 26308 22428 26314
rect 22376 26250 22428 26256
rect 22388 26042 22416 26250
rect 22376 26036 22428 26042
rect 22376 25978 22428 25984
rect 22622 25596 22930 25605
rect 22622 25594 22628 25596
rect 22684 25594 22708 25596
rect 22764 25594 22788 25596
rect 22844 25594 22868 25596
rect 22924 25594 22930 25596
rect 22684 25542 22686 25594
rect 22866 25542 22868 25594
rect 22622 25540 22628 25542
rect 22684 25540 22708 25542
rect 22764 25540 22788 25542
rect 22844 25540 22868 25542
rect 22924 25540 22930 25542
rect 22622 25531 22930 25540
rect 22284 25424 22336 25430
rect 22284 25366 22336 25372
rect 21916 25288 21968 25294
rect 21916 25230 21968 25236
rect 21824 24948 21876 24954
rect 21824 24890 21876 24896
rect 21836 24274 21864 24890
rect 21928 24750 21956 25230
rect 22008 25152 22060 25158
rect 22008 25094 22060 25100
rect 22020 24954 22048 25094
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 22008 24812 22060 24818
rect 22008 24754 22060 24760
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21824 24268 21876 24274
rect 21824 24210 21876 24216
rect 21836 23526 21864 24210
rect 21928 23730 21956 24550
rect 22020 24342 22048 24754
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 22020 23730 22048 24278
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 21916 23724 21968 23730
rect 21916 23666 21968 23672
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 21824 23520 21876 23526
rect 21824 23462 21876 23468
rect 21824 22568 21876 22574
rect 21824 22510 21876 22516
rect 21836 22234 21864 22510
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 22112 22094 22140 24142
rect 22204 23322 22232 24618
rect 22296 24274 22324 25366
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22296 22642 22324 24210
rect 22388 23254 22416 24890
rect 22622 24508 22930 24517
rect 22622 24506 22628 24508
rect 22684 24506 22708 24508
rect 22764 24506 22788 24508
rect 22844 24506 22868 24508
rect 22924 24506 22930 24508
rect 22684 24454 22686 24506
rect 22866 24454 22868 24506
rect 22622 24452 22628 24454
rect 22684 24452 22708 24454
rect 22764 24452 22788 24454
rect 22844 24452 22868 24454
rect 22924 24452 22930 24454
rect 22622 24443 22930 24452
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22480 23866 22508 24006
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 22622 23420 22930 23429
rect 22622 23418 22628 23420
rect 22684 23418 22708 23420
rect 22764 23418 22788 23420
rect 22844 23418 22868 23420
rect 22924 23418 22930 23420
rect 22684 23366 22686 23418
rect 22866 23366 22868 23418
rect 22622 23364 22628 23366
rect 22684 23364 22708 23366
rect 22764 23364 22788 23366
rect 22844 23364 22868 23366
rect 22924 23364 22930 23366
rect 22622 23355 22930 23364
rect 22376 23248 22428 23254
rect 22376 23190 22428 23196
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22622 22332 22930 22341
rect 22622 22330 22628 22332
rect 22684 22330 22708 22332
rect 22764 22330 22788 22332
rect 22844 22330 22868 22332
rect 22924 22330 22930 22332
rect 22684 22278 22686 22330
rect 22866 22278 22868 22330
rect 22622 22276 22628 22278
rect 22684 22276 22708 22278
rect 22764 22276 22788 22278
rect 22844 22276 22868 22278
rect 22924 22276 22930 22278
rect 22622 22267 22930 22276
rect 22112 22066 22232 22094
rect 22098 21992 22154 22001
rect 21824 21956 21876 21962
rect 22098 21927 22154 21936
rect 21824 21898 21876 21904
rect 21836 21865 21864 21898
rect 21822 21856 21878 21865
rect 21822 21791 21878 21800
rect 21836 21078 21864 21791
rect 22112 21146 22140 21927
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 21824 21072 21876 21078
rect 22204 21026 22232 22066
rect 22468 22024 22520 22030
rect 22744 22024 22796 22030
rect 22468 21966 22520 21972
rect 22742 21992 22744 22001
rect 22796 21992 22798 22001
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 21824 21014 21876 21020
rect 22112 20998 22232 21026
rect 22112 18426 22140 20998
rect 22296 20942 22324 21490
rect 22480 21350 22508 21966
rect 22742 21927 22798 21936
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22622 21244 22930 21253
rect 22622 21242 22628 21244
rect 22684 21242 22708 21244
rect 22764 21242 22788 21244
rect 22844 21242 22868 21244
rect 22924 21242 22930 21244
rect 22684 21190 22686 21242
rect 22866 21190 22868 21242
rect 22622 21188 22628 21190
rect 22684 21188 22708 21190
rect 22764 21188 22788 21190
rect 22844 21188 22868 21190
rect 22924 21188 22930 21190
rect 22622 21179 22930 21188
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22204 20466 22232 20878
rect 23032 20534 23060 26794
rect 23400 26518 23428 26930
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 23112 26240 23164 26246
rect 23112 26182 23164 26188
rect 23020 20528 23072 20534
rect 23020 20470 23072 20476
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22622 20156 22930 20165
rect 22622 20154 22628 20156
rect 22684 20154 22708 20156
rect 22764 20154 22788 20156
rect 22844 20154 22868 20156
rect 22924 20154 22930 20156
rect 22684 20102 22686 20154
rect 22866 20102 22868 20154
rect 22622 20100 22628 20102
rect 22684 20100 22708 20102
rect 22764 20100 22788 20102
rect 22844 20100 22868 20102
rect 22924 20100 22930 20102
rect 22190 20088 22246 20097
rect 22622 20091 22930 20100
rect 22190 20023 22246 20032
rect 22376 20052 22428 20058
rect 22204 19990 22232 20023
rect 22376 19994 22428 20000
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 22284 19780 22336 19786
rect 22284 19722 22336 19728
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22190 18320 22246 18329
rect 22100 18284 22152 18290
rect 22190 18255 22246 18264
rect 22100 18226 22152 18232
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21836 17377 21864 18090
rect 21822 17368 21878 17377
rect 21822 17303 21878 17312
rect 21836 17202 21864 17303
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21824 15088 21876 15094
rect 21824 15030 21876 15036
rect 21836 12238 21864 15030
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21928 14346 21956 14894
rect 22008 14408 22060 14414
rect 22006 14376 22008 14385
rect 22060 14376 22062 14385
rect 21916 14340 21968 14346
rect 22006 14311 22062 14320
rect 21916 14282 21968 14288
rect 22112 13326 22140 18226
rect 22204 15094 22232 18255
rect 22296 17490 22324 19722
rect 22388 19378 22416 19994
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22388 18329 22416 18770
rect 22480 18766 22508 19790
rect 23032 19786 23060 20470
rect 23020 19780 23072 19786
rect 23020 19722 23072 19728
rect 22622 19068 22930 19077
rect 22622 19066 22628 19068
rect 22684 19066 22708 19068
rect 22764 19066 22788 19068
rect 22844 19066 22868 19068
rect 22924 19066 22930 19068
rect 22684 19014 22686 19066
rect 22866 19014 22868 19066
rect 22622 19012 22628 19014
rect 22684 19012 22708 19014
rect 22764 19012 22788 19014
rect 22844 19012 22868 19014
rect 22924 19012 22930 19014
rect 22622 19003 22930 19012
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22374 18320 22430 18329
rect 22374 18255 22430 18264
rect 22480 18086 22508 18702
rect 22468 18080 22520 18086
rect 22374 18048 22430 18057
rect 22468 18022 22520 18028
rect 22374 17983 22430 17992
rect 22388 17678 22416 17983
rect 22622 17980 22930 17989
rect 22622 17978 22628 17980
rect 22684 17978 22708 17980
rect 22764 17978 22788 17980
rect 22844 17978 22868 17980
rect 22924 17978 22930 17980
rect 22684 17926 22686 17978
rect 22866 17926 22868 17978
rect 22622 17924 22628 17926
rect 22684 17924 22708 17926
rect 22764 17924 22788 17926
rect 22844 17924 22868 17926
rect 22924 17924 22930 17926
rect 22622 17915 22930 17924
rect 22928 17876 22980 17882
rect 22928 17818 22980 17824
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 22376 17672 22428 17678
rect 22428 17620 22508 17626
rect 22376 17614 22508 17620
rect 22388 17598 22508 17614
rect 22296 17462 22416 17490
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22296 16522 22324 16934
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22284 16108 22336 16114
rect 22388 16096 22416 17462
rect 22336 16068 22416 16096
rect 22284 16050 22336 16056
rect 22296 15434 22324 16050
rect 22284 15428 22336 15434
rect 22284 15370 22336 15376
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22480 14464 22508 17598
rect 22940 17270 22968 17818
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 22622 16892 22930 16901
rect 22622 16890 22628 16892
rect 22684 16890 22708 16892
rect 22764 16890 22788 16892
rect 22844 16890 22868 16892
rect 22924 16890 22930 16892
rect 22684 16838 22686 16890
rect 22866 16838 22868 16890
rect 22622 16836 22628 16838
rect 22684 16836 22708 16838
rect 22764 16836 22788 16838
rect 22844 16836 22868 16838
rect 22924 16836 22930 16838
rect 22622 16827 22930 16836
rect 23032 16794 23060 17818
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 22622 15804 22930 15813
rect 22622 15802 22628 15804
rect 22684 15802 22708 15804
rect 22764 15802 22788 15804
rect 22844 15802 22868 15804
rect 22924 15802 22930 15804
rect 22684 15750 22686 15802
rect 22866 15750 22868 15802
rect 22622 15748 22628 15750
rect 22684 15748 22708 15750
rect 22764 15748 22788 15750
rect 22844 15748 22868 15750
rect 22924 15748 22930 15750
rect 22622 15739 22930 15748
rect 23032 15502 23060 16730
rect 23124 16250 23152 26182
rect 23400 25974 23428 26454
rect 24228 26450 24256 26726
rect 24216 26444 24268 26450
rect 24216 26386 24268 26392
rect 23848 26240 23900 26246
rect 23848 26182 23900 26188
rect 23388 25968 23440 25974
rect 23388 25910 23440 25916
rect 23860 25906 23888 26182
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23940 25220 23992 25226
rect 23940 25162 23992 25168
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23216 24206 23244 25094
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 23400 24410 23428 24686
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23400 23594 23428 24346
rect 23768 24206 23796 24550
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23860 24138 23888 24550
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 23216 22234 23244 22374
rect 23204 22228 23256 22234
rect 23204 22170 23256 22176
rect 23296 21548 23348 21554
rect 23400 21536 23428 23530
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23584 23186 23612 23462
rect 23572 23180 23624 23186
rect 23572 23122 23624 23128
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23492 22710 23520 22986
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23480 22704 23532 22710
rect 23480 22646 23532 22652
rect 23584 22166 23612 22918
rect 23860 22794 23888 24074
rect 23952 23254 23980 25162
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 24136 23526 24164 24210
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 23940 23248 23992 23254
rect 23940 23190 23992 23196
rect 23768 22766 23888 22794
rect 23664 22636 23716 22642
rect 23768 22624 23796 22766
rect 23716 22596 23796 22624
rect 23664 22578 23716 22584
rect 23768 22438 23796 22596
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23756 22432 23808 22438
rect 23756 22374 23808 22380
rect 23572 22160 23624 22166
rect 23572 22102 23624 22108
rect 23860 21962 23888 22578
rect 23952 22574 23980 23190
rect 24136 22794 24164 23462
rect 24136 22778 24256 22794
rect 24136 22772 24268 22778
rect 24136 22766 24216 22772
rect 24216 22714 24268 22720
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 23952 22137 23980 22510
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 24044 22166 24072 22374
rect 24032 22160 24084 22166
rect 23938 22128 23994 22137
rect 24032 22102 24084 22108
rect 23938 22063 23994 22072
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23348 21508 23428 21536
rect 23296 21490 23348 21496
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23676 21146 23704 21422
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23860 21078 23888 21898
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23860 20262 23888 20878
rect 24136 20602 24164 22578
rect 24216 22500 24268 22506
rect 24216 22442 24268 22448
rect 24228 21962 24256 22442
rect 24216 21956 24268 21962
rect 24216 21898 24268 21904
rect 24320 20641 24348 32710
rect 24412 32230 24440 33254
rect 24400 32224 24452 32230
rect 24400 32166 24452 32172
rect 27160 29572 27212 29578
rect 27160 29514 27212 29520
rect 26424 29504 26476 29510
rect 26424 29446 26476 29452
rect 26436 29238 26464 29446
rect 26424 29232 26476 29238
rect 26424 29174 26476 29180
rect 26792 29164 26844 29170
rect 26792 29106 26844 29112
rect 26804 28558 26832 29106
rect 27172 28762 27200 29514
rect 27160 28756 27212 28762
rect 27160 28698 27212 28704
rect 26792 28552 26844 28558
rect 26792 28494 26844 28500
rect 27356 26382 27384 33254
rect 33612 33114 33640 33458
rect 36268 33380 36320 33386
rect 36268 33322 36320 33328
rect 35900 33312 35952 33318
rect 35900 33254 35952 33260
rect 35912 33130 35940 33254
rect 33600 33108 33652 33114
rect 33600 33050 33652 33056
rect 35820 33102 35940 33130
rect 35820 32910 35848 33102
rect 35808 32904 35860 32910
rect 35808 32846 35860 32852
rect 36280 32892 36308 33322
rect 37740 33312 37792 33318
rect 37740 33254 37792 33260
rect 37070 33212 37378 33221
rect 37070 33210 37076 33212
rect 37132 33210 37156 33212
rect 37212 33210 37236 33212
rect 37292 33210 37316 33212
rect 37372 33210 37378 33212
rect 37132 33158 37134 33210
rect 37314 33158 37316 33210
rect 37070 33156 37076 33158
rect 37132 33156 37156 33158
rect 37212 33156 37236 33158
rect 37292 33156 37316 33158
rect 37372 33156 37378 33158
rect 37070 33147 37378 33156
rect 37752 32910 37780 33254
rect 38948 33114 38976 33458
rect 38936 33108 38988 33114
rect 38936 33050 38988 33056
rect 36452 32904 36504 32910
rect 36280 32864 36452 32892
rect 32956 32768 33008 32774
rect 32956 32710 33008 32716
rect 35716 32768 35768 32774
rect 35716 32710 35768 32716
rect 29846 32668 30154 32677
rect 29846 32666 29852 32668
rect 29908 32666 29932 32668
rect 29988 32666 30012 32668
rect 30068 32666 30092 32668
rect 30148 32666 30154 32668
rect 29908 32614 29910 32666
rect 30090 32614 30092 32666
rect 29846 32612 29852 32614
rect 29908 32612 29932 32614
rect 29988 32612 30012 32614
rect 30068 32612 30092 32614
rect 30148 32612 30154 32614
rect 29846 32603 30154 32612
rect 29846 31580 30154 31589
rect 29846 31578 29852 31580
rect 29908 31578 29932 31580
rect 29988 31578 30012 31580
rect 30068 31578 30092 31580
rect 30148 31578 30154 31580
rect 29908 31526 29910 31578
rect 30090 31526 30092 31578
rect 29846 31524 29852 31526
rect 29908 31524 29932 31526
rect 29988 31524 30012 31526
rect 30068 31524 30092 31526
rect 30148 31524 30154 31526
rect 29846 31515 30154 31524
rect 29846 30492 30154 30501
rect 29846 30490 29852 30492
rect 29908 30490 29932 30492
rect 29988 30490 30012 30492
rect 30068 30490 30092 30492
rect 30148 30490 30154 30492
rect 29908 30438 29910 30490
rect 30090 30438 30092 30490
rect 29846 30436 29852 30438
rect 29908 30436 29932 30438
rect 29988 30436 30012 30438
rect 30068 30436 30092 30438
rect 30148 30436 30154 30438
rect 29846 30427 30154 30436
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27540 29102 27568 29650
rect 30196 29504 30248 29510
rect 30196 29446 30248 29452
rect 29846 29404 30154 29413
rect 29846 29402 29852 29404
rect 29908 29402 29932 29404
rect 29988 29402 30012 29404
rect 30068 29402 30092 29404
rect 30148 29402 30154 29404
rect 29908 29350 29910 29402
rect 30090 29350 30092 29402
rect 29846 29348 29852 29350
rect 29908 29348 29932 29350
rect 29988 29348 30012 29350
rect 30068 29348 30092 29350
rect 30148 29348 30154 29350
rect 29846 29339 30154 29348
rect 27528 29096 27580 29102
rect 27528 29038 27580 29044
rect 28908 29096 28960 29102
rect 28908 29038 28960 29044
rect 27436 28960 27488 28966
rect 27436 28902 27488 28908
rect 27448 28762 27476 28902
rect 27436 28756 27488 28762
rect 27436 28698 27488 28704
rect 27540 28558 27568 29038
rect 27528 28552 27580 28558
rect 27528 28494 27580 28500
rect 27344 26376 27396 26382
rect 27344 26318 27396 26324
rect 28724 25900 28776 25906
rect 28724 25842 28776 25848
rect 27436 25696 27488 25702
rect 27436 25638 27488 25644
rect 26330 25392 26386 25401
rect 26330 25327 26332 25336
rect 26384 25327 26386 25336
rect 26332 25298 26384 25304
rect 26608 25220 26660 25226
rect 26608 25162 26660 25168
rect 26620 24954 26648 25162
rect 26608 24948 26660 24954
rect 26608 24890 26660 24896
rect 24490 24848 24546 24857
rect 24490 24783 24492 24792
rect 24544 24783 24546 24792
rect 25044 24812 25096 24818
rect 24492 24754 24544 24760
rect 25044 24754 25096 24760
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 24768 24064 24820 24070
rect 24768 24006 24820 24012
rect 24584 23792 24636 23798
rect 24584 23734 24636 23740
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 24412 22386 24440 23666
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24504 23089 24532 23598
rect 24596 23118 24624 23734
rect 24676 23520 24728 23526
rect 24676 23462 24728 23468
rect 24584 23112 24636 23118
rect 24490 23080 24546 23089
rect 24584 23054 24636 23060
rect 24490 23015 24492 23024
rect 24544 23015 24546 23024
rect 24492 22986 24544 22992
rect 24504 22955 24532 22986
rect 24688 22778 24716 23462
rect 24780 23100 24808 24006
rect 24952 23112 25004 23118
rect 24780 23072 24952 23100
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24596 22522 24624 22714
rect 24676 22636 24728 22642
rect 24780 22624 24808 23072
rect 24952 23054 25004 23060
rect 24728 22596 24808 22624
rect 24952 22636 25004 22642
rect 24676 22578 24728 22584
rect 24952 22578 25004 22584
rect 24596 22494 24808 22522
rect 24964 22506 24992 22578
rect 24412 22358 24624 22386
rect 24596 22234 24624 22358
rect 24584 22228 24636 22234
rect 24584 22170 24636 22176
rect 24490 22128 24546 22137
rect 24490 22063 24546 22072
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24412 21146 24440 21966
rect 24504 21894 24532 22063
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24504 21593 24532 21830
rect 24490 21584 24546 21593
rect 24490 21519 24546 21528
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 24306 20632 24362 20641
rect 24124 20596 24176 20602
rect 24306 20567 24362 20576
rect 24124 20538 24176 20544
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23308 18442 23336 20198
rect 23756 19712 23808 19718
rect 23400 19638 23612 19666
rect 23756 19654 23808 19660
rect 23400 19514 23428 19638
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 23308 18414 23428 18442
rect 23294 17232 23350 17241
rect 23294 17167 23296 17176
rect 23348 17167 23350 17176
rect 23296 17138 23348 17144
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23216 16182 23244 16934
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 23400 15178 23428 18414
rect 23492 16590 23520 19450
rect 23584 18834 23612 19638
rect 23768 19242 23796 19654
rect 23756 19236 23808 19242
rect 23756 19178 23808 19184
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23584 17882 23612 18770
rect 23768 18766 23796 19178
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23848 17604 23900 17610
rect 23848 17546 23900 17552
rect 23480 16584 23532 16590
rect 23480 16526 23532 16532
rect 23860 15706 23888 17546
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23216 15150 23428 15178
rect 22622 14716 22930 14725
rect 22622 14714 22628 14716
rect 22684 14714 22708 14716
rect 22764 14714 22788 14716
rect 22844 14714 22868 14716
rect 22924 14714 22930 14716
rect 22684 14662 22686 14714
rect 22866 14662 22868 14714
rect 22622 14660 22628 14662
rect 22684 14660 22708 14662
rect 22764 14660 22788 14662
rect 22844 14660 22868 14662
rect 22924 14660 22930 14662
rect 22622 14651 22930 14660
rect 22296 14436 22508 14464
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22204 13172 22232 14214
rect 22112 13144 22232 13172
rect 22112 12850 22140 13144
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22296 12345 22324 14436
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22388 13462 22416 14282
rect 23020 14272 23072 14278
rect 23020 14214 23072 14220
rect 22836 14068 22888 14074
rect 23032 14056 23060 14214
rect 22888 14028 23060 14056
rect 22836 14010 22888 14016
rect 22622 13628 22930 13637
rect 22622 13626 22628 13628
rect 22684 13626 22708 13628
rect 22764 13626 22788 13628
rect 22844 13626 22868 13628
rect 22924 13626 22930 13628
rect 22684 13574 22686 13626
rect 22866 13574 22868 13626
rect 22622 13572 22628 13574
rect 22684 13572 22708 13574
rect 22764 13572 22788 13574
rect 22844 13572 22868 13574
rect 22924 13572 22930 13574
rect 22622 13563 22930 13572
rect 22376 13456 22428 13462
rect 22376 13398 22428 13404
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 22480 12986 22508 13398
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 23032 12782 23060 14028
rect 23216 13870 23244 15150
rect 23492 14414 23520 15370
rect 24044 15026 24072 15438
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23584 14618 23612 14894
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 22622 12540 22930 12549
rect 22622 12538 22628 12540
rect 22684 12538 22708 12540
rect 22764 12538 22788 12540
rect 22844 12538 22868 12540
rect 22924 12538 22930 12540
rect 22684 12486 22686 12538
rect 22866 12486 22868 12538
rect 22622 12484 22628 12486
rect 22684 12484 22708 12486
rect 22764 12484 22788 12486
rect 22844 12484 22868 12486
rect 22924 12484 22930 12486
rect 22622 12475 22930 12484
rect 22282 12336 22338 12345
rect 22282 12271 22338 12280
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 23216 12170 23244 12922
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 23204 12164 23256 12170
rect 23204 12106 23256 12112
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 21928 10810 21956 10950
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 21928 10674 21956 10746
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 22112 10062 22140 12106
rect 23478 11792 23534 11801
rect 23478 11727 23480 11736
rect 23532 11727 23534 11736
rect 23480 11698 23532 11704
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 22388 10742 22416 11018
rect 22376 10736 22428 10742
rect 22376 10678 22428 10684
rect 22100 10056 22152 10062
rect 21914 10024 21970 10033
rect 22100 9998 22152 10004
rect 21914 9959 21970 9968
rect 21928 9722 21956 9959
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22480 9654 22508 11630
rect 22622 11452 22930 11461
rect 22622 11450 22628 11452
rect 22684 11450 22708 11452
rect 22764 11450 22788 11452
rect 22844 11450 22868 11452
rect 22924 11450 22930 11452
rect 22684 11398 22686 11450
rect 22866 11398 22868 11450
rect 22622 11396 22628 11398
rect 22684 11396 22708 11398
rect 22764 11396 22788 11398
rect 22844 11396 22868 11398
rect 22924 11396 22930 11398
rect 22622 11387 22930 11396
rect 23584 10606 23612 14554
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 23952 14074 23980 14418
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 24044 13530 24072 14962
rect 24136 13870 24164 20538
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 24228 18766 24256 19110
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24412 15910 24440 18566
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24688 17814 24716 18158
rect 24676 17808 24728 17814
rect 24676 17750 24728 17756
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24688 16574 24716 16730
rect 24596 16546 24716 16574
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24412 15586 24440 15846
rect 24504 15706 24532 16118
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24308 15564 24360 15570
rect 24412 15558 24532 15586
rect 24308 15506 24360 15512
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24228 12918 24256 14758
rect 24320 13308 24348 15506
rect 24400 14000 24452 14006
rect 24400 13942 24452 13948
rect 24412 13530 24440 13942
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24400 13320 24452 13326
rect 24320 13280 24400 13308
rect 24400 13262 24452 13268
rect 24504 13274 24532 15558
rect 24596 15502 24624 16546
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24688 16182 24716 16390
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24596 13394 24624 15438
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24688 15094 24716 15302
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 24780 14618 24808 22494
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24872 21554 24900 21830
rect 24964 21690 24992 21966
rect 25056 21729 25084 24754
rect 25320 24744 25372 24750
rect 25320 24686 25372 24692
rect 25136 24336 25188 24342
rect 25136 24278 25188 24284
rect 25148 24070 25176 24278
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25148 23866 25176 24006
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25226 23080 25282 23089
rect 25226 23015 25282 23024
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 25148 22642 25176 22918
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 25042 21720 25098 21729
rect 24952 21684 25004 21690
rect 25042 21655 25098 21664
rect 24952 21626 25004 21632
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24964 21486 24992 21626
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24964 21146 24992 21286
rect 24952 21140 25004 21146
rect 24952 21082 25004 21088
rect 25240 20942 25268 23015
rect 25332 22778 25360 24686
rect 26436 24410 26464 24754
rect 26792 24608 26844 24614
rect 26792 24550 26844 24556
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25516 23225 25544 23598
rect 26056 23520 26108 23526
rect 26056 23462 26108 23468
rect 25502 23216 25558 23225
rect 25502 23151 25558 23160
rect 25596 23180 25648 23186
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 25516 22642 25544 23151
rect 25596 23122 25648 23128
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25608 22574 25636 23122
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25780 23112 25832 23118
rect 25780 23054 25832 23060
rect 25700 22778 25728 23054
rect 25792 22982 25820 23054
rect 25780 22976 25832 22982
rect 25780 22918 25832 22924
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25700 22166 25728 22714
rect 25792 22506 25820 22918
rect 25780 22500 25832 22506
rect 25780 22442 25832 22448
rect 25688 22160 25740 22166
rect 25688 22102 25740 22108
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25504 21888 25556 21894
rect 25504 21830 25556 21836
rect 25516 21622 25544 21830
rect 25608 21690 25636 21966
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25504 21616 25556 21622
rect 25504 21558 25556 21564
rect 25228 20936 25280 20942
rect 25228 20878 25280 20884
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25700 20534 25728 20742
rect 25688 20528 25740 20534
rect 25688 20470 25740 20476
rect 25688 20256 25740 20262
rect 25056 20182 25268 20210
rect 25688 20198 25740 20204
rect 25056 20058 25084 20182
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24872 19802 24900 19858
rect 24872 19774 25084 19802
rect 25148 19786 25176 19994
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24872 18426 24900 19314
rect 25056 19310 25084 19774
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25148 19446 25176 19722
rect 25136 19440 25188 19446
rect 25136 19382 25188 19388
rect 25044 19304 25096 19310
rect 25044 19246 25096 19252
rect 25056 18426 25084 19246
rect 24860 18420 24912 18426
rect 24860 18362 24912 18368
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 24872 17202 24900 18362
rect 24952 18352 25004 18358
rect 24952 18294 25004 18300
rect 24964 17882 24992 18294
rect 25240 18222 25268 20182
rect 25700 19922 25728 20198
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25792 18766 25820 22034
rect 26068 22030 26096 23462
rect 26252 22642 26280 24006
rect 26436 23730 26464 24210
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26436 22642 26464 23054
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26424 22636 26476 22642
rect 26424 22578 26476 22584
rect 26240 22500 26292 22506
rect 26240 22442 26292 22448
rect 26056 22024 26108 22030
rect 26056 21966 26108 21972
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 25872 21412 25924 21418
rect 25872 21354 25924 21360
rect 25884 20346 25912 21354
rect 25976 20466 26004 21898
rect 26068 21622 26096 21966
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26160 21729 26188 21830
rect 26146 21720 26202 21729
rect 26146 21655 26202 21664
rect 26056 21616 26108 21622
rect 26056 21558 26108 21564
rect 26160 21078 26188 21655
rect 26252 21554 26280 22442
rect 26528 22030 26556 24142
rect 26804 24138 26832 24550
rect 27448 24177 27476 25638
rect 28736 25294 28764 25842
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 28080 25152 28132 25158
rect 28080 25094 28132 25100
rect 28092 24818 28120 25094
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 27988 24404 28040 24410
rect 27988 24346 28040 24352
rect 27434 24168 27490 24177
rect 26792 24132 26844 24138
rect 27434 24103 27490 24112
rect 26792 24074 26844 24080
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26608 23588 26660 23594
rect 26608 23530 26660 23536
rect 26620 23118 26648 23530
rect 26988 23118 27016 23666
rect 27448 23322 27476 24103
rect 28000 23730 28028 24346
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 28092 23662 28120 24754
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 28368 24138 28396 24550
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28356 24132 28408 24138
rect 28356 24074 28408 24080
rect 28080 23656 28132 23662
rect 28080 23598 28132 23604
rect 27528 23588 27580 23594
rect 27528 23530 27580 23536
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 26608 23112 26660 23118
rect 26884 23112 26936 23118
rect 26608 23054 26660 23060
rect 26882 23080 26884 23089
rect 26976 23112 27028 23118
rect 26936 23080 26938 23089
rect 26976 23054 27028 23060
rect 26882 23015 26938 23024
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 26516 22024 26568 22030
rect 26516 21966 26568 21972
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 26884 21616 26936 21622
rect 26884 21558 26936 21564
rect 27066 21584 27122 21593
rect 26240 21548 26292 21554
rect 26240 21490 26292 21496
rect 26896 21418 26924 21558
rect 27172 21554 27200 21966
rect 27356 21894 27384 22510
rect 27540 22094 27568 23530
rect 28736 23526 28764 24210
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 27620 23316 27672 23322
rect 27620 23258 27672 23264
rect 27448 22066 27568 22094
rect 27344 21888 27396 21894
rect 27344 21830 27396 21836
rect 27066 21519 27122 21528
rect 27160 21548 27212 21554
rect 27080 21486 27108 21519
rect 27160 21490 27212 21496
rect 27252 21548 27304 21554
rect 27252 21490 27304 21496
rect 27068 21480 27120 21486
rect 27068 21422 27120 21428
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 26884 21412 26936 21418
rect 26884 21354 26936 21360
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26148 21072 26200 21078
rect 26148 21014 26200 21020
rect 26252 20942 26280 21286
rect 26528 21078 26556 21354
rect 27172 21162 27200 21490
rect 27080 21146 27200 21162
rect 27264 21146 27292 21490
rect 27356 21418 27384 21830
rect 27344 21412 27396 21418
rect 27344 21354 27396 21360
rect 27068 21140 27200 21146
rect 27120 21134 27200 21140
rect 27252 21140 27304 21146
rect 27068 21082 27120 21088
rect 27252 21082 27304 21088
rect 26516 21072 26568 21078
rect 26516 21014 26568 21020
rect 27356 21010 27384 21354
rect 27344 21004 27396 21010
rect 27344 20946 27396 20952
rect 27448 20942 27476 22066
rect 27632 21622 27660 23258
rect 28080 23248 28132 23254
rect 28080 23190 28132 23196
rect 27988 23044 28040 23050
rect 27988 22986 28040 22992
rect 28000 22710 28028 22986
rect 27988 22704 28040 22710
rect 27988 22646 28040 22652
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27816 22166 27844 22374
rect 27804 22160 27856 22166
rect 27804 22102 27856 22108
rect 28000 22094 28028 22646
rect 27908 22066 28028 22094
rect 27908 21690 27936 22066
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 27804 21684 27856 21690
rect 27804 21626 27856 21632
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27620 21616 27672 21622
rect 27620 21558 27672 21564
rect 27540 21418 27568 21558
rect 27528 21412 27580 21418
rect 27528 21354 27580 21360
rect 27816 21350 27844 21626
rect 27896 21548 27948 21554
rect 27896 21490 27948 21496
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 26148 20596 26200 20602
rect 26148 20538 26200 20544
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 26160 20346 26188 20538
rect 25884 20318 26188 20346
rect 25884 19854 25912 20318
rect 26252 19854 26280 20878
rect 27448 20262 27476 20878
rect 27632 20466 27660 21286
rect 27908 21078 27936 21490
rect 28000 21146 28028 21966
rect 28092 21486 28120 23190
rect 28632 23180 28684 23186
rect 28632 23122 28684 23128
rect 28172 23112 28224 23118
rect 28172 23054 28224 23060
rect 28184 22012 28212 23054
rect 28540 22976 28592 22982
rect 28540 22918 28592 22924
rect 28552 22234 28580 22918
rect 28644 22642 28672 23122
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28540 22228 28592 22234
rect 28540 22170 28592 22176
rect 28264 22024 28316 22030
rect 28184 21984 28264 22012
rect 28184 21554 28212 21984
rect 28264 21966 28316 21972
rect 28356 21956 28408 21962
rect 28356 21898 28408 21904
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 28080 21480 28132 21486
rect 28080 21422 28132 21428
rect 27988 21140 28040 21146
rect 27988 21082 28040 21088
rect 27896 21072 27948 21078
rect 27896 21014 27948 21020
rect 28262 20632 28318 20641
rect 28368 20602 28396 21898
rect 28736 20942 28764 23462
rect 28816 22976 28868 22982
rect 28816 22918 28868 22924
rect 28828 22166 28856 22918
rect 28816 22160 28868 22166
rect 28816 22102 28868 22108
rect 28816 21344 28868 21350
rect 28816 21286 28868 21292
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28262 20567 28318 20576
rect 28356 20596 28408 20602
rect 28276 20534 28304 20567
rect 28356 20538 28408 20544
rect 27896 20528 27948 20534
rect 27896 20470 27948 20476
rect 28264 20528 28316 20534
rect 28264 20470 28316 20476
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 27908 19990 27936 20470
rect 28080 20460 28132 20466
rect 28080 20402 28132 20408
rect 27620 19984 27672 19990
rect 27620 19926 27672 19932
rect 27896 19984 27948 19990
rect 27896 19926 27948 19932
rect 25872 19848 25924 19854
rect 25872 19790 25924 19796
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 27344 19712 27396 19718
rect 27250 19680 27306 19689
rect 27344 19654 27396 19660
rect 27250 19615 27306 19624
rect 27264 19446 27292 19615
rect 27252 19440 27304 19446
rect 27252 19382 27304 19388
rect 26608 19236 26660 19242
rect 26608 19178 26660 19184
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 25688 18352 25740 18358
rect 25688 18294 25740 18300
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 25700 17338 25728 18294
rect 25976 17678 26004 18702
rect 26068 18358 26096 18906
rect 26160 18698 26188 19110
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26056 18352 26108 18358
rect 26056 18294 26108 18300
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 26160 17678 26188 18158
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 25964 17672 26016 17678
rect 25964 17614 26016 17620
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 23768 12442 23796 12854
rect 23848 12640 23900 12646
rect 23848 12582 23900 12588
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23768 11830 23796 12038
rect 23860 11898 23888 12582
rect 24412 12306 24440 13262
rect 24504 13246 24716 13274
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23848 11212 23900 11218
rect 23848 11154 23900 11160
rect 23860 11082 23888 11154
rect 24412 11150 24440 12038
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 22622 10364 22930 10373
rect 22622 10362 22628 10364
rect 22684 10362 22708 10364
rect 22764 10362 22788 10364
rect 22844 10362 22868 10364
rect 22924 10362 22930 10364
rect 22684 10310 22686 10362
rect 22866 10310 22868 10362
rect 22622 10308 22628 10310
rect 22684 10308 22708 10310
rect 22764 10308 22788 10310
rect 22844 10308 22868 10310
rect 22924 10308 22930 10310
rect 22622 10299 22930 10308
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 23860 9586 23888 11018
rect 24504 10742 24532 11630
rect 24492 10736 24544 10742
rect 24492 10678 24544 10684
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24504 10146 24532 10542
rect 24596 10266 24624 12242
rect 24688 11218 24716 13246
rect 24780 11898 24808 13806
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24964 11150 24992 17070
rect 25056 16998 25084 17274
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25792 16674 25820 16730
rect 25976 16726 26004 17614
rect 25424 16658 25820 16674
rect 25964 16720 26016 16726
rect 25964 16662 26016 16668
rect 25412 16652 25820 16658
rect 25464 16646 25820 16652
rect 25412 16594 25464 16600
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 25424 14346 25452 15846
rect 26252 15706 26280 18090
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 26240 15700 26292 15706
rect 26240 15642 26292 15648
rect 25964 14816 26016 14822
rect 25964 14758 26016 14764
rect 25412 14340 25464 14346
rect 25412 14282 25464 14288
rect 25976 13258 26004 14758
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26252 13326 26280 13874
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 25412 13184 25464 13190
rect 25412 13126 25464 13132
rect 25424 12170 25452 13126
rect 26148 12232 26200 12238
rect 26146 12200 26148 12209
rect 26200 12200 26202 12209
rect 25412 12164 25464 12170
rect 26146 12135 26202 12144
rect 25412 12106 25464 12112
rect 26160 11898 26188 12135
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 25504 11076 25556 11082
rect 25504 11018 25556 11024
rect 25516 10674 25544 11018
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24504 10118 24716 10146
rect 26252 10130 26280 13262
rect 26436 12238 26464 16934
rect 26620 16574 26648 19178
rect 26792 18624 26844 18630
rect 26792 18566 26844 18572
rect 26804 17105 26832 18566
rect 27356 18329 27384 19654
rect 27632 18698 27660 19926
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27804 19780 27856 19786
rect 27804 19722 27856 19728
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 27342 18320 27398 18329
rect 27342 18255 27398 18264
rect 27436 18284 27488 18290
rect 27436 18226 27488 18232
rect 27344 17604 27396 17610
rect 27448 17592 27476 18226
rect 27724 18222 27752 19654
rect 27816 19514 27844 19722
rect 27804 19508 27856 19514
rect 27804 19450 27856 19456
rect 27908 19394 27936 19790
rect 27816 19366 27936 19394
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27396 17564 27476 17592
rect 27344 17546 27396 17552
rect 26790 17096 26846 17105
rect 26790 17031 26846 17040
rect 26976 16992 27028 16998
rect 26976 16934 27028 16940
rect 26528 16546 26648 16574
rect 26528 12986 26556 16546
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26620 15366 26648 16050
rect 26608 15360 26660 15366
rect 26660 15308 26832 15314
rect 26608 15302 26832 15308
rect 26620 15286 26832 15302
rect 26804 14414 26832 15286
rect 26988 15162 27016 16934
rect 27356 15978 27384 17546
rect 27712 16584 27764 16590
rect 27816 16574 27844 19366
rect 28092 18970 28120 20402
rect 28276 19854 28304 20470
rect 28828 19854 28856 21286
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28080 18964 28132 18970
rect 28080 18906 28132 18912
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 27816 16546 27936 16574
rect 27712 16526 27764 16532
rect 27620 16448 27672 16454
rect 27620 16390 27672 16396
rect 27632 16114 27660 16390
rect 27620 16108 27672 16114
rect 27620 16050 27672 16056
rect 27344 15972 27396 15978
rect 27344 15914 27396 15920
rect 27528 15972 27580 15978
rect 27528 15914 27580 15920
rect 27540 15502 27568 15914
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 26976 15156 27028 15162
rect 26976 15098 27028 15104
rect 26988 14890 27016 15098
rect 26976 14884 27028 14890
rect 26976 14826 27028 14832
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 26792 14408 26844 14414
rect 26792 14350 26844 14356
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26712 14006 26740 14214
rect 26700 14000 26752 14006
rect 26700 13942 26752 13948
rect 26804 13530 26832 14350
rect 27068 13864 27120 13870
rect 27068 13806 27120 13812
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26516 12980 26568 12986
rect 26516 12922 26568 12928
rect 26882 12336 26938 12345
rect 26882 12271 26938 12280
rect 26896 12238 26924 12271
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 27080 11830 27108 13806
rect 27068 11824 27120 11830
rect 27068 11766 27120 11772
rect 27356 11354 27384 14554
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27448 14074 27476 14350
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27540 13870 27568 15438
rect 27632 15026 27660 16050
rect 27724 16046 27752 16526
rect 27712 16040 27764 16046
rect 27712 15982 27764 15988
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27724 14906 27752 15982
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27632 14878 27752 14906
rect 27632 14550 27660 14878
rect 27620 14544 27672 14550
rect 27620 14486 27672 14492
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27632 14113 27660 14350
rect 27618 14104 27674 14113
rect 27618 14039 27674 14048
rect 27816 13938 27844 15030
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27620 12640 27672 12646
rect 27620 12582 27672 12588
rect 27632 12102 27660 12582
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 26516 11008 26568 11014
rect 26516 10950 26568 10956
rect 26528 10130 26556 10950
rect 27160 10600 27212 10606
rect 27160 10542 27212 10548
rect 27172 10130 27200 10542
rect 27712 10192 27764 10198
rect 27712 10134 27764 10140
rect 24688 9994 24716 10118
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 27160 10124 27212 10130
rect 27160 10066 27212 10072
rect 24676 9988 24728 9994
rect 24676 9930 24728 9936
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 24688 9518 24716 9930
rect 26424 9920 26476 9926
rect 26424 9862 26476 9868
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 22622 9276 22930 9285
rect 22622 9274 22628 9276
rect 22684 9274 22708 9276
rect 22764 9274 22788 9276
rect 22844 9274 22868 9276
rect 22924 9274 22930 9276
rect 22684 9222 22686 9274
rect 22866 9222 22868 9274
rect 22622 9220 22628 9222
rect 22684 9220 22708 9222
rect 22764 9220 22788 9222
rect 22844 9220 22868 9222
rect 22924 9220 22930 9222
rect 22622 9211 22930 9220
rect 26436 8974 26464 9862
rect 27252 9376 27304 9382
rect 27252 9318 27304 9324
rect 27264 9110 27292 9318
rect 27252 9104 27304 9110
rect 27252 9046 27304 9052
rect 27264 8974 27292 9046
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 26436 8634 26464 8910
rect 26424 8628 26476 8634
rect 26424 8570 26476 8576
rect 22622 8188 22930 8197
rect 22622 8186 22628 8188
rect 22684 8186 22708 8188
rect 22764 8186 22788 8188
rect 22844 8186 22868 8188
rect 22924 8186 22930 8188
rect 22684 8134 22686 8186
rect 22866 8134 22868 8186
rect 22622 8132 22628 8134
rect 22684 8132 22708 8134
rect 22764 8132 22788 8134
rect 22844 8132 22868 8134
rect 22924 8132 22930 8134
rect 22622 8123 22930 8132
rect 26436 8090 26464 8570
rect 27724 8294 27752 10134
rect 27712 8288 27764 8294
rect 27712 8230 27764 8236
rect 26424 8084 26476 8090
rect 26424 8026 26476 8032
rect 27816 7954 27844 11630
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 27802 7848 27858 7857
rect 27802 7783 27804 7792
rect 27856 7783 27858 7792
rect 27804 7754 27856 7760
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 22622 7100 22930 7109
rect 22622 7098 22628 7100
rect 22684 7098 22708 7100
rect 22764 7098 22788 7100
rect 22844 7098 22868 7100
rect 22924 7098 22930 7100
rect 22684 7046 22686 7098
rect 22866 7046 22868 7098
rect 22622 7044 22628 7046
rect 22684 7044 22708 7046
rect 22764 7044 22788 7046
rect 22844 7044 22868 7046
rect 22924 7044 22930 7046
rect 22622 7035 22930 7044
rect 27632 6866 27660 7482
rect 27712 7336 27764 7342
rect 27712 7278 27764 7284
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27724 6662 27752 7278
rect 27816 6798 27844 7754
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27712 6656 27764 6662
rect 27712 6598 27764 6604
rect 25964 6248 26016 6254
rect 25964 6190 26016 6196
rect 22622 6012 22930 6021
rect 22622 6010 22628 6012
rect 22684 6010 22708 6012
rect 22764 6010 22788 6012
rect 22844 6010 22868 6012
rect 22924 6010 22930 6012
rect 22684 5958 22686 6010
rect 22866 5958 22868 6010
rect 22622 5956 22628 5958
rect 22684 5956 22708 5958
rect 22764 5956 22788 5958
rect 22844 5956 22868 5958
rect 22924 5956 22930 5958
rect 22622 5947 22930 5956
rect 25976 5914 26004 6190
rect 27724 6186 27752 6598
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 27712 6180 27764 6186
rect 27712 6122 27764 6128
rect 27816 5914 27844 6326
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 27804 5908 27856 5914
rect 27804 5850 27856 5856
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26252 5370 26280 5646
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 26240 5364 26292 5370
rect 26240 5306 26292 5312
rect 19720 3058 19748 5306
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 24768 5092 24820 5098
rect 24768 5034 24820 5040
rect 22622 4924 22930 4933
rect 22622 4922 22628 4924
rect 22684 4922 22708 4924
rect 22764 4922 22788 4924
rect 22844 4922 22868 4924
rect 22924 4922 22930 4924
rect 22684 4870 22686 4922
rect 22866 4870 22868 4922
rect 22622 4868 22628 4870
rect 22684 4868 22708 4870
rect 22764 4868 22788 4870
rect 22844 4868 22868 4870
rect 22924 4868 22930 4870
rect 22622 4859 22930 4868
rect 24780 4826 24808 5034
rect 24860 5024 24912 5030
rect 24860 4966 24912 4972
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24872 4622 24900 4966
rect 25884 4826 25912 5170
rect 25872 4820 25924 4826
rect 25872 4762 25924 4768
rect 26332 4752 26384 4758
rect 26332 4694 26384 4700
rect 24860 4616 24912 4622
rect 24858 4584 24860 4593
rect 24912 4584 24914 4593
rect 26344 4554 26372 4694
rect 24858 4519 24914 4528
rect 25412 4548 25464 4554
rect 25412 4490 25464 4496
rect 26332 4548 26384 4554
rect 26332 4490 26384 4496
rect 25320 4072 25372 4078
rect 25320 4014 25372 4020
rect 25332 3942 25360 4014
rect 25424 4010 25452 4490
rect 25412 4004 25464 4010
rect 25412 3946 25464 3952
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 22622 3836 22930 3845
rect 22622 3834 22628 3836
rect 22684 3834 22708 3836
rect 22764 3834 22788 3836
rect 22844 3834 22868 3836
rect 22924 3834 22930 3836
rect 22684 3782 22686 3834
rect 22866 3782 22868 3834
rect 22622 3780 22628 3782
rect 22684 3780 22708 3782
rect 22764 3780 22788 3782
rect 22844 3780 22868 3782
rect 22924 3780 22930 3782
rect 22622 3771 22930 3780
rect 23124 3602 23152 3878
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 25332 3534 25360 3878
rect 26344 3738 26372 4490
rect 26988 4282 27016 5170
rect 27160 4480 27212 4486
rect 27160 4422 27212 4428
rect 27252 4480 27304 4486
rect 27252 4422 27304 4428
rect 26976 4276 27028 4282
rect 26976 4218 27028 4224
rect 27172 4146 27200 4422
rect 27264 4214 27292 4422
rect 27252 4208 27304 4214
rect 27252 4150 27304 4156
rect 27160 4140 27212 4146
rect 27160 4082 27212 4088
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 27264 3466 27292 4150
rect 27252 3460 27304 3466
rect 27252 3402 27304 3408
rect 27908 3058 27936 16546
rect 28000 15434 28028 18634
rect 28092 18222 28120 18906
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28080 18216 28132 18222
rect 28080 18158 28132 18164
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 28092 16182 28120 17138
rect 28184 16590 28212 18226
rect 28724 17740 28776 17746
rect 28724 17682 28776 17688
rect 28354 17368 28410 17377
rect 28354 17303 28410 17312
rect 28368 17202 28396 17303
rect 28356 17196 28408 17202
rect 28356 17138 28408 17144
rect 28172 16584 28224 16590
rect 28172 16526 28224 16532
rect 28632 16448 28684 16454
rect 28632 16390 28684 16396
rect 28080 16176 28132 16182
rect 28080 16118 28132 16124
rect 27988 15428 28040 15434
rect 27988 15370 28040 15376
rect 28644 15094 28672 16390
rect 28632 15088 28684 15094
rect 28632 15030 28684 15036
rect 28080 14816 28132 14822
rect 28080 14758 28132 14764
rect 28092 14482 28120 14758
rect 28080 14476 28132 14482
rect 28080 14418 28132 14424
rect 28448 14272 28500 14278
rect 28448 14214 28500 14220
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 28092 13530 28120 13806
rect 28080 13524 28132 13530
rect 28080 13466 28132 13472
rect 28264 12096 28316 12102
rect 28264 12038 28316 12044
rect 28276 11830 28304 12038
rect 28264 11824 28316 11830
rect 28264 11766 28316 11772
rect 28172 11076 28224 11082
rect 28172 11018 28224 11024
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 27988 9444 28040 9450
rect 27988 9386 28040 9392
rect 28000 7274 28028 9386
rect 28092 7886 28120 9454
rect 28184 9382 28212 11018
rect 28264 10192 28316 10198
rect 28264 10134 28316 10140
rect 28172 9376 28224 9382
rect 28172 9318 28224 9324
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 28184 8566 28212 8910
rect 28172 8560 28224 8566
rect 28172 8502 28224 8508
rect 28276 8378 28304 10134
rect 28460 9654 28488 14214
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 28644 11354 28672 12242
rect 28632 11348 28684 11354
rect 28632 11290 28684 11296
rect 28736 10130 28764 17682
rect 28816 17060 28868 17066
rect 28816 17002 28868 17008
rect 28828 16454 28856 17002
rect 28816 16448 28868 16454
rect 28816 16390 28868 16396
rect 28828 15366 28856 16390
rect 28816 15360 28868 15366
rect 28816 15302 28868 15308
rect 28828 15065 28856 15302
rect 28814 15056 28870 15065
rect 28814 14991 28870 15000
rect 28724 10124 28776 10130
rect 28724 10066 28776 10072
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28448 9648 28500 9654
rect 28448 9590 28500 9596
rect 28736 8906 28764 9930
rect 28724 8900 28776 8906
rect 28724 8842 28776 8848
rect 28736 8634 28764 8842
rect 28724 8628 28776 8634
rect 28724 8570 28776 8576
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 28184 8350 28304 8378
rect 28184 8090 28212 8350
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28092 7546 28120 7822
rect 28080 7540 28132 7546
rect 28080 7482 28132 7488
rect 28184 7290 28212 8026
rect 28460 7750 28488 8434
rect 28816 8288 28868 8294
rect 28816 8230 28868 8236
rect 28632 7948 28684 7954
rect 28632 7890 28684 7896
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28262 7440 28318 7449
rect 28262 7375 28264 7384
rect 28316 7375 28318 7384
rect 28264 7346 28316 7352
rect 28460 7342 28488 7686
rect 28644 7410 28672 7890
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 28736 7546 28764 7822
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28632 7404 28684 7410
rect 28632 7346 28684 7352
rect 28356 7336 28408 7342
rect 27988 7268 28040 7274
rect 28184 7262 28304 7290
rect 28356 7278 28408 7284
rect 28448 7336 28500 7342
rect 28448 7278 28500 7284
rect 27988 7210 28040 7216
rect 28000 6934 28028 7210
rect 28080 7200 28132 7206
rect 28080 7142 28132 7148
rect 27988 6928 28040 6934
rect 27988 6870 28040 6876
rect 28092 6322 28120 7142
rect 28276 6662 28304 7262
rect 28368 6730 28396 7278
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 28264 6656 28316 6662
rect 28264 6598 28316 6604
rect 28276 6390 28304 6598
rect 28264 6384 28316 6390
rect 28264 6326 28316 6332
rect 28080 6316 28132 6322
rect 28080 6258 28132 6264
rect 28092 3602 28120 6258
rect 28644 5710 28672 7346
rect 28828 7041 28856 8230
rect 28814 7032 28870 7041
rect 28814 6967 28870 6976
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 28736 5778 28764 6054
rect 28920 5914 28948 29038
rect 29846 28316 30154 28325
rect 29846 28314 29852 28316
rect 29908 28314 29932 28316
rect 29988 28314 30012 28316
rect 30068 28314 30092 28316
rect 30148 28314 30154 28316
rect 29908 28262 29910 28314
rect 30090 28262 30092 28314
rect 29846 28260 29852 28262
rect 29908 28260 29932 28262
rect 29988 28260 30012 28262
rect 30068 28260 30092 28262
rect 30148 28260 30154 28262
rect 29846 28251 30154 28260
rect 29846 27228 30154 27237
rect 29846 27226 29852 27228
rect 29908 27226 29932 27228
rect 29988 27226 30012 27228
rect 30068 27226 30092 27228
rect 30148 27226 30154 27228
rect 29908 27174 29910 27226
rect 30090 27174 30092 27226
rect 29846 27172 29852 27174
rect 29908 27172 29932 27174
rect 29988 27172 30012 27174
rect 30068 27172 30092 27174
rect 30148 27172 30154 27174
rect 29846 27163 30154 27172
rect 29846 26140 30154 26149
rect 29846 26138 29852 26140
rect 29908 26138 29932 26140
rect 29988 26138 30012 26140
rect 30068 26138 30092 26140
rect 30148 26138 30154 26140
rect 29908 26086 29910 26138
rect 30090 26086 30092 26138
rect 29846 26084 29852 26086
rect 29908 26084 29932 26086
rect 29988 26084 30012 26086
rect 30068 26084 30092 26086
rect 30148 26084 30154 26086
rect 29846 26075 30154 26084
rect 29552 25288 29604 25294
rect 29552 25230 29604 25236
rect 29564 24886 29592 25230
rect 29846 25052 30154 25061
rect 29846 25050 29852 25052
rect 29908 25050 29932 25052
rect 29988 25050 30012 25052
rect 30068 25050 30092 25052
rect 30148 25050 30154 25052
rect 29908 24998 29910 25050
rect 30090 24998 30092 25050
rect 29846 24996 29852 24998
rect 29908 24996 29932 24998
rect 29988 24996 30012 24998
rect 30068 24996 30092 24998
rect 30148 24996 30154 24998
rect 29846 24987 30154 24996
rect 29552 24880 29604 24886
rect 29552 24822 29604 24828
rect 29000 24812 29052 24818
rect 29000 24754 29052 24760
rect 29012 24410 29040 24754
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 30012 24608 30064 24614
rect 30012 24550 30064 24556
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29460 24064 29512 24070
rect 29460 24006 29512 24012
rect 29472 23662 29500 24006
rect 29564 23730 29592 24142
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29748 23712 29776 24550
rect 30024 24410 30052 24550
rect 30012 24404 30064 24410
rect 30012 24346 30064 24352
rect 29846 23964 30154 23973
rect 29846 23962 29852 23964
rect 29908 23962 29932 23964
rect 29988 23962 30012 23964
rect 30068 23962 30092 23964
rect 30148 23962 30154 23964
rect 29908 23910 29910 23962
rect 30090 23910 30092 23962
rect 29846 23908 29852 23910
rect 29908 23908 29932 23910
rect 29988 23908 30012 23910
rect 30068 23908 30092 23910
rect 30148 23908 30154 23910
rect 29846 23899 30154 23908
rect 29828 23724 29880 23730
rect 29748 23684 29828 23712
rect 29276 23656 29328 23662
rect 29276 23598 29328 23604
rect 29460 23656 29512 23662
rect 29460 23598 29512 23604
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 29012 22030 29040 23054
rect 29092 22432 29144 22438
rect 29092 22374 29144 22380
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 29012 21078 29040 21966
rect 29000 21072 29052 21078
rect 29000 21014 29052 21020
rect 29104 20806 29132 22374
rect 29288 21010 29316 23598
rect 29656 22438 29684 23598
rect 29644 22432 29696 22438
rect 29644 22374 29696 22380
rect 29748 22098 29776 23684
rect 29828 23666 29880 23672
rect 29846 22876 30154 22885
rect 29846 22874 29852 22876
rect 29908 22874 29932 22876
rect 29988 22874 30012 22876
rect 30068 22874 30092 22876
rect 30148 22874 30154 22876
rect 29908 22822 29910 22874
rect 30090 22822 30092 22874
rect 29846 22820 29852 22822
rect 29908 22820 29932 22822
rect 29988 22820 30012 22822
rect 30068 22820 30092 22822
rect 30148 22820 30154 22822
rect 29846 22811 30154 22820
rect 30104 22568 30156 22574
rect 30104 22510 30156 22516
rect 30116 22234 30144 22510
rect 30104 22228 30156 22234
rect 30104 22170 30156 22176
rect 29736 22092 29788 22098
rect 29736 22034 29788 22040
rect 29460 21888 29512 21894
rect 29460 21830 29512 21836
rect 29366 21448 29422 21457
rect 29366 21383 29368 21392
rect 29420 21383 29422 21392
rect 29368 21354 29420 21360
rect 29276 21004 29328 21010
rect 29276 20946 29328 20952
rect 29092 20800 29144 20806
rect 29092 20742 29144 20748
rect 29472 20602 29500 21830
rect 29748 20874 29776 22034
rect 29846 21788 30154 21797
rect 29846 21786 29852 21788
rect 29908 21786 29932 21788
rect 29988 21786 30012 21788
rect 30068 21786 30092 21788
rect 30148 21786 30154 21788
rect 29908 21734 29910 21786
rect 30090 21734 30092 21786
rect 29846 21732 29852 21734
rect 29908 21732 29932 21734
rect 29988 21732 30012 21734
rect 30068 21732 30092 21734
rect 30148 21732 30154 21734
rect 29846 21723 30154 21732
rect 30208 21622 30236 29446
rect 30288 27328 30340 27334
rect 30288 27270 30340 27276
rect 30300 26790 30328 27270
rect 30288 26784 30340 26790
rect 30288 26726 30340 26732
rect 30300 25974 30328 26726
rect 30288 25968 30340 25974
rect 30288 25910 30340 25916
rect 30932 25696 30984 25702
rect 30932 25638 30984 25644
rect 30944 25294 30972 25638
rect 30932 25288 30984 25294
rect 30932 25230 30984 25236
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 31312 24750 31340 25094
rect 31772 24818 31800 25230
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31300 24744 31352 24750
rect 31300 24686 31352 24692
rect 31772 24410 31800 24754
rect 31852 24676 31904 24682
rect 31852 24618 31904 24624
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 31208 24132 31260 24138
rect 31208 24074 31260 24080
rect 31220 23866 31248 24074
rect 31760 24064 31812 24070
rect 31760 24006 31812 24012
rect 31208 23860 31260 23866
rect 31208 23802 31260 23808
rect 31392 23044 31444 23050
rect 31392 22986 31444 22992
rect 31404 22778 31432 22986
rect 31392 22772 31444 22778
rect 31392 22714 31444 22720
rect 31576 22432 31628 22438
rect 31576 22374 31628 22380
rect 31588 22098 31616 22374
rect 31576 22092 31628 22098
rect 31576 22034 31628 22040
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 30196 21616 30248 21622
rect 30196 21558 30248 21564
rect 29828 21344 29880 21350
rect 29828 21286 29880 21292
rect 29840 21010 29868 21286
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 29736 20868 29788 20874
rect 29736 20810 29788 20816
rect 29846 20700 30154 20709
rect 29846 20698 29852 20700
rect 29908 20698 29932 20700
rect 29988 20698 30012 20700
rect 30068 20698 30092 20700
rect 30148 20698 30154 20700
rect 29908 20646 29910 20698
rect 30090 20646 30092 20698
rect 29846 20644 29852 20646
rect 29908 20644 29932 20646
rect 29988 20644 30012 20646
rect 30068 20644 30092 20646
rect 30148 20644 30154 20646
rect 29846 20635 30154 20644
rect 29460 20596 29512 20602
rect 29460 20538 29512 20544
rect 30104 20528 30156 20534
rect 30104 20470 30156 20476
rect 30116 20058 30144 20470
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 29000 19780 29052 19786
rect 29000 19722 29052 19728
rect 29012 18970 29040 19722
rect 29846 19612 30154 19621
rect 29846 19610 29852 19612
rect 29908 19610 29932 19612
rect 29988 19610 30012 19612
rect 30068 19610 30092 19612
rect 30148 19610 30154 19612
rect 29908 19558 29910 19610
rect 30090 19558 30092 19610
rect 29846 19556 29852 19558
rect 29908 19556 29932 19558
rect 29988 19556 30012 19558
rect 30068 19556 30092 19558
rect 30148 19556 30154 19558
rect 29846 19547 30154 19556
rect 30208 19310 30236 21558
rect 30484 21486 30512 21966
rect 31300 21956 31352 21962
rect 31300 21898 31352 21904
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 30472 21480 30524 21486
rect 30472 21422 30524 21428
rect 30484 19854 30512 21422
rect 30576 20874 30604 21830
rect 31312 21146 31340 21898
rect 31588 21554 31616 22034
rect 31576 21548 31628 21554
rect 31576 21490 31628 21496
rect 31300 21140 31352 21146
rect 31300 21082 31352 21088
rect 31772 21010 31800 24006
rect 31864 23730 31892 24618
rect 31852 23724 31904 23730
rect 31852 23666 31904 23672
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 31864 23186 31892 23666
rect 32128 23520 32180 23526
rect 32128 23462 32180 23468
rect 31852 23180 31904 23186
rect 31852 23122 31904 23128
rect 32140 23050 32168 23462
rect 32692 23050 32720 23666
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 32680 23044 32732 23050
rect 32680 22986 32732 22992
rect 32692 22642 32720 22986
rect 32864 22976 32916 22982
rect 32864 22918 32916 22924
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 31864 21418 31892 22578
rect 32312 21888 32364 21894
rect 32312 21830 32364 21836
rect 31852 21412 31904 21418
rect 31852 21354 31904 21360
rect 32036 21344 32088 21350
rect 32036 21286 32088 21292
rect 32048 21010 32076 21286
rect 31760 21004 31812 21010
rect 31760 20946 31812 20952
rect 32036 21004 32088 21010
rect 32036 20946 32088 20952
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 31024 20392 31076 20398
rect 31024 20334 31076 20340
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30656 19848 30708 19854
rect 30656 19790 30708 19796
rect 30564 19440 30616 19446
rect 30564 19382 30616 19388
rect 29460 19304 29512 19310
rect 29460 19246 29512 19252
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 29472 18834 29500 19246
rect 29460 18828 29512 18834
rect 29460 18770 29512 18776
rect 29644 18624 29696 18630
rect 29644 18566 29696 18572
rect 29656 18426 29684 18566
rect 29846 18524 30154 18533
rect 29846 18522 29852 18524
rect 29908 18522 29932 18524
rect 29988 18522 30012 18524
rect 30068 18522 30092 18524
rect 30148 18522 30154 18524
rect 29908 18470 29910 18522
rect 30090 18470 30092 18522
rect 29846 18468 29852 18470
rect 29908 18468 29932 18470
rect 29988 18468 30012 18470
rect 30068 18468 30092 18470
rect 30148 18468 30154 18470
rect 29846 18459 30154 18468
rect 30208 18426 30236 19246
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 29644 18420 29696 18426
rect 29644 18362 29696 18368
rect 30196 18420 30248 18426
rect 30196 18362 30248 18368
rect 29276 18216 29328 18222
rect 29276 18158 29328 18164
rect 29288 17134 29316 18158
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29276 17128 29328 17134
rect 29276 17070 29328 17076
rect 28998 15464 29054 15473
rect 29054 15434 29132 15450
rect 29054 15428 29144 15434
rect 29054 15422 29092 15428
rect 28998 15399 29054 15408
rect 29012 14618 29040 15399
rect 29092 15370 29144 15376
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 29104 13954 29132 14894
rect 29012 13926 29132 13954
rect 29012 11694 29040 13926
rect 29092 13796 29144 13802
rect 29092 13738 29144 13744
rect 29104 12374 29132 13738
rect 29092 12368 29144 12374
rect 29092 12310 29144 12316
rect 29000 11688 29052 11694
rect 29000 11630 29052 11636
rect 29196 10742 29224 17070
rect 29644 17060 29696 17066
rect 29644 17002 29696 17008
rect 29552 16652 29604 16658
rect 29552 16594 29604 16600
rect 29564 16289 29592 16594
rect 29550 16280 29606 16289
rect 29550 16215 29606 16224
rect 29276 16040 29328 16046
rect 29656 16017 29684 17002
rect 29748 16590 29776 17478
rect 29846 17436 30154 17445
rect 29846 17434 29852 17436
rect 29908 17434 29932 17436
rect 29988 17434 30012 17436
rect 30068 17434 30092 17436
rect 30148 17434 30154 17436
rect 29908 17382 29910 17434
rect 30090 17382 30092 17434
rect 29846 17380 29852 17382
rect 29908 17380 29932 17382
rect 29988 17380 30012 17382
rect 30068 17380 30092 17382
rect 30148 17380 30154 17382
rect 29846 17371 30154 17380
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 30116 16794 30144 17070
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 29736 16584 29788 16590
rect 30392 16574 30420 19110
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 30484 18290 30512 18702
rect 30472 18284 30524 18290
rect 30472 18226 30524 18232
rect 30576 17814 30604 19382
rect 30668 18358 30696 19790
rect 31036 19514 31064 20334
rect 31208 19780 31260 19786
rect 31208 19722 31260 19728
rect 31944 19780 31996 19786
rect 31944 19722 31996 19728
rect 31116 19712 31168 19718
rect 31116 19654 31168 19660
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 31024 19372 31076 19378
rect 31024 19314 31076 19320
rect 30656 18352 30708 18358
rect 30656 18294 30708 18300
rect 30932 18284 30984 18290
rect 30932 18226 30984 18232
rect 30564 17808 30616 17814
rect 30564 17750 30616 17756
rect 30392 16546 30512 16574
rect 29736 16526 29788 16532
rect 29748 16250 29776 16526
rect 29846 16348 30154 16357
rect 29846 16346 29852 16348
rect 29908 16346 29932 16348
rect 29988 16346 30012 16348
rect 30068 16346 30092 16348
rect 30148 16346 30154 16348
rect 29908 16294 29910 16346
rect 30090 16294 30092 16346
rect 29846 16292 29852 16294
rect 29908 16292 29932 16294
rect 29988 16292 30012 16294
rect 30068 16292 30092 16294
rect 30148 16292 30154 16294
rect 29846 16283 30154 16292
rect 29736 16244 29788 16250
rect 29736 16186 29788 16192
rect 29276 15982 29328 15988
rect 29642 16008 29698 16017
rect 29092 10736 29144 10742
rect 29092 10678 29144 10684
rect 29184 10736 29236 10742
rect 29184 10678 29236 10684
rect 29104 7750 29132 10678
rect 29288 9654 29316 15982
rect 29642 15943 29698 15952
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 29460 15564 29512 15570
rect 29460 15506 29512 15512
rect 29472 13326 29500 15506
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29460 13320 29512 13326
rect 29460 13262 29512 13268
rect 29472 12918 29500 13262
rect 29460 12912 29512 12918
rect 29460 12854 29512 12860
rect 29564 12306 29592 15438
rect 29846 15260 30154 15269
rect 29846 15258 29852 15260
rect 29908 15258 29932 15260
rect 29988 15258 30012 15260
rect 30068 15258 30092 15260
rect 30148 15258 30154 15260
rect 29908 15206 29910 15258
rect 30090 15206 30092 15258
rect 29846 15204 29852 15206
rect 29908 15204 29932 15206
rect 29988 15204 30012 15206
rect 30068 15204 30092 15206
rect 30148 15204 30154 15206
rect 29846 15195 30154 15204
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29748 14074 29776 14350
rect 29846 14172 30154 14181
rect 29846 14170 29852 14172
rect 29908 14170 29932 14172
rect 29988 14170 30012 14172
rect 30068 14170 30092 14172
rect 30148 14170 30154 14172
rect 29908 14118 29910 14170
rect 30090 14118 30092 14170
rect 29846 14116 29852 14118
rect 29908 14116 29932 14118
rect 29988 14116 30012 14118
rect 30068 14116 30092 14118
rect 30148 14116 30154 14118
rect 29846 14107 30154 14116
rect 29736 14068 29788 14074
rect 29736 14010 29788 14016
rect 29644 14000 29696 14006
rect 29644 13942 29696 13948
rect 29656 13530 29684 13942
rect 30392 13818 30420 15846
rect 30484 15162 30512 16546
rect 30944 16114 30972 18226
rect 31036 17082 31064 19314
rect 31128 18290 31156 19654
rect 31220 18290 31248 19722
rect 31392 18760 31444 18766
rect 31392 18702 31444 18708
rect 31116 18284 31168 18290
rect 31116 18226 31168 18232
rect 31208 18284 31260 18290
rect 31208 18226 31260 18232
rect 31206 17640 31262 17649
rect 31206 17575 31208 17584
rect 31260 17575 31262 17584
rect 31208 17546 31260 17552
rect 31404 17202 31432 18702
rect 31956 18358 31984 19722
rect 32036 18692 32088 18698
rect 32036 18634 32088 18640
rect 31944 18352 31996 18358
rect 31944 18294 31996 18300
rect 31576 17808 31628 17814
rect 31576 17750 31628 17756
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31036 17054 31432 17082
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 31036 16590 31064 16934
rect 31312 16658 31340 16934
rect 31300 16652 31352 16658
rect 31300 16594 31352 16600
rect 31024 16584 31076 16590
rect 31024 16526 31076 16532
rect 30932 16108 30984 16114
rect 30932 16050 30984 16056
rect 30564 16040 30616 16046
rect 30564 15982 30616 15988
rect 30472 15156 30524 15162
rect 30472 15098 30524 15104
rect 30484 14482 30512 15098
rect 30576 15094 30604 15982
rect 31036 15722 31064 16526
rect 30944 15694 31064 15722
rect 30564 15088 30616 15094
rect 30564 15030 30616 15036
rect 30472 14476 30524 14482
rect 30472 14418 30524 14424
rect 30944 13977 30972 15694
rect 31404 15586 31432 17054
rect 31312 15558 31432 15586
rect 30930 13968 30986 13977
rect 30930 13903 30986 13912
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 31208 13932 31260 13938
rect 31208 13874 31260 13880
rect 30208 13790 30420 13818
rect 30748 13864 30800 13870
rect 30748 13806 30800 13812
rect 31036 13818 31064 13874
rect 30208 13734 30236 13790
rect 30196 13728 30248 13734
rect 30196 13670 30248 13676
rect 30380 13728 30432 13734
rect 30380 13670 30432 13676
rect 29644 13524 29696 13530
rect 29644 13466 29696 13472
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 29846 13084 30154 13093
rect 29846 13082 29852 13084
rect 29908 13082 29932 13084
rect 29988 13082 30012 13084
rect 30068 13082 30092 13084
rect 30148 13082 30154 13084
rect 29908 13030 29910 13082
rect 30090 13030 30092 13082
rect 29846 13028 29852 13030
rect 29908 13028 29932 13030
rect 29988 13028 30012 13030
rect 30068 13028 30092 13030
rect 30148 13028 30154 13030
rect 29846 13019 30154 13028
rect 30300 12986 30328 13262
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 29828 12912 29880 12918
rect 29826 12880 29828 12889
rect 29880 12880 29882 12889
rect 29826 12815 29882 12824
rect 30392 12442 30420 13670
rect 30760 13394 30788 13806
rect 31036 13790 31156 13818
rect 30748 13388 30800 13394
rect 30748 13330 30800 13336
rect 30380 12436 30432 12442
rect 30380 12378 30432 12384
rect 30656 12436 30708 12442
rect 30656 12378 30708 12384
rect 30288 12368 30340 12374
rect 30288 12310 30340 12316
rect 29552 12300 29604 12306
rect 29552 12242 29604 12248
rect 29564 11830 29592 12242
rect 29846 11996 30154 12005
rect 29846 11994 29852 11996
rect 29908 11994 29932 11996
rect 29988 11994 30012 11996
rect 30068 11994 30092 11996
rect 30148 11994 30154 11996
rect 29908 11942 29910 11994
rect 30090 11942 30092 11994
rect 29846 11940 29852 11942
rect 29908 11940 29932 11942
rect 29988 11940 30012 11942
rect 30068 11940 30092 11942
rect 30148 11940 30154 11942
rect 29846 11931 30154 11940
rect 29552 11824 29604 11830
rect 29552 11766 29604 11772
rect 30104 11824 30156 11830
rect 30104 11766 30156 11772
rect 30116 11082 30144 11766
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30104 11076 30156 11082
rect 30104 11018 30156 11024
rect 29846 10908 30154 10917
rect 29846 10906 29852 10908
rect 29908 10906 29932 10908
rect 29988 10906 30012 10908
rect 30068 10906 30092 10908
rect 30148 10906 30154 10908
rect 29908 10854 29910 10906
rect 30090 10854 30092 10906
rect 29846 10852 29852 10854
rect 29908 10852 29932 10854
rect 29988 10852 30012 10854
rect 30068 10852 30092 10854
rect 30148 10852 30154 10854
rect 29846 10843 30154 10852
rect 30208 10606 30236 11630
rect 30300 11218 30328 12310
rect 30668 12238 30696 12378
rect 30656 12232 30708 12238
rect 30656 12174 30708 12180
rect 30668 11898 30696 12174
rect 30656 11892 30708 11898
rect 30656 11834 30708 11840
rect 30760 11778 30788 13330
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30852 11898 30880 13262
rect 31024 13252 31076 13258
rect 30944 13212 31024 13240
rect 30944 12646 30972 13212
rect 31024 13194 31076 13200
rect 31128 12986 31156 13790
rect 31116 12980 31168 12986
rect 31116 12922 31168 12928
rect 30932 12640 30984 12646
rect 30932 12582 30984 12588
rect 31024 12164 31076 12170
rect 31024 12106 31076 12112
rect 30840 11892 30892 11898
rect 30840 11834 30892 11840
rect 30564 11756 30616 11762
rect 30760 11750 30880 11778
rect 30564 11698 30616 11704
rect 30378 11656 30434 11665
rect 30378 11591 30434 11600
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 30392 11150 30420 11591
rect 30576 11286 30604 11698
rect 30564 11280 30616 11286
rect 30564 11222 30616 11228
rect 30380 11144 30432 11150
rect 30380 11086 30432 11092
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 30196 10600 30248 10606
rect 30196 10542 30248 10548
rect 29368 10192 29420 10198
rect 29368 10134 29420 10140
rect 29276 9648 29328 9654
rect 29276 9590 29328 9596
rect 29380 9042 29408 10134
rect 29368 9036 29420 9042
rect 29368 8978 29420 8984
rect 29380 8634 29408 8978
rect 29368 8628 29420 8634
rect 29368 8570 29420 8576
rect 29564 8344 29592 10542
rect 30380 10532 30432 10538
rect 30380 10474 30432 10480
rect 30286 9888 30342 9897
rect 29846 9820 30154 9829
rect 30286 9823 30342 9832
rect 29846 9818 29852 9820
rect 29908 9818 29932 9820
rect 29988 9818 30012 9820
rect 30068 9818 30092 9820
rect 30148 9818 30154 9820
rect 29908 9766 29910 9818
rect 30090 9766 30092 9818
rect 29846 9764 29852 9766
rect 29908 9764 29932 9766
rect 29988 9764 30012 9766
rect 30068 9764 30092 9766
rect 30148 9764 30154 9766
rect 29846 9755 30154 9764
rect 30196 9376 30248 9382
rect 30196 9318 30248 9324
rect 29734 9072 29790 9081
rect 29644 9036 29696 9042
rect 29734 9007 29790 9016
rect 29644 8978 29696 8984
rect 29656 8634 29684 8978
rect 29748 8974 29776 9007
rect 29736 8968 29788 8974
rect 29736 8910 29788 8916
rect 29846 8732 30154 8741
rect 29846 8730 29852 8732
rect 29908 8730 29932 8732
rect 29988 8730 30012 8732
rect 30068 8730 30092 8732
rect 30148 8730 30154 8732
rect 29908 8678 29910 8730
rect 30090 8678 30092 8730
rect 29846 8676 29852 8678
rect 29908 8676 29932 8678
rect 29988 8676 30012 8678
rect 30068 8676 30092 8678
rect 30148 8676 30154 8678
rect 29846 8667 30154 8676
rect 29644 8628 29696 8634
rect 29644 8570 29696 8576
rect 29644 8356 29696 8362
rect 29564 8316 29644 8344
rect 29644 8298 29696 8304
rect 29460 7948 29512 7954
rect 29460 7890 29512 7896
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 29184 7472 29236 7478
rect 29184 7414 29236 7420
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 29104 6798 29132 7142
rect 29092 6792 29144 6798
rect 29092 6734 29144 6740
rect 29196 6662 29224 7414
rect 29472 6866 29500 7890
rect 29656 7410 29684 8298
rect 29736 7880 29788 7886
rect 29736 7822 29788 7828
rect 29748 7546 29776 7822
rect 29846 7644 30154 7653
rect 29846 7642 29852 7644
rect 29908 7642 29932 7644
rect 29988 7642 30012 7644
rect 30068 7642 30092 7644
rect 30148 7642 30154 7644
rect 29908 7590 29910 7642
rect 30090 7590 30092 7642
rect 29846 7588 29852 7590
rect 29908 7588 29932 7590
rect 29988 7588 30012 7590
rect 30068 7588 30092 7590
rect 30148 7588 30154 7590
rect 29846 7579 30154 7588
rect 29736 7540 29788 7546
rect 29736 7482 29788 7488
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29656 7206 29684 7346
rect 29644 7200 29696 7206
rect 29644 7142 29696 7148
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 29184 6656 29236 6662
rect 29184 6598 29236 6604
rect 29368 6656 29420 6662
rect 29368 6598 29420 6604
rect 29380 6322 29408 6598
rect 29368 6316 29420 6322
rect 29368 6258 29420 6264
rect 29472 6254 29500 6802
rect 29460 6248 29512 6254
rect 29460 6190 29512 6196
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 28632 5704 28684 5710
rect 28632 5646 28684 5652
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 29196 5166 29224 5510
rect 29656 5234 29684 7142
rect 30208 6798 30236 9318
rect 30300 8498 30328 9823
rect 30392 9382 30420 10474
rect 30472 10260 30524 10266
rect 30472 10202 30524 10208
rect 30484 10169 30512 10202
rect 30470 10160 30526 10169
rect 30470 10095 30526 10104
rect 30472 10056 30524 10062
rect 30576 10044 30604 11222
rect 30748 10600 30800 10606
rect 30748 10542 30800 10548
rect 30656 10532 30708 10538
rect 30656 10474 30708 10480
rect 30668 10266 30696 10474
rect 30656 10260 30708 10266
rect 30656 10202 30708 10208
rect 30524 10016 30604 10044
rect 30472 9998 30524 10004
rect 30380 9376 30432 9382
rect 30380 9318 30432 9324
rect 30484 9042 30512 9998
rect 30656 9716 30708 9722
rect 30760 9704 30788 10542
rect 30852 10130 30880 11750
rect 30930 11656 30986 11665
rect 30930 11591 30932 11600
rect 30984 11591 30986 11600
rect 30932 11562 30984 11568
rect 30944 11354 30972 11562
rect 30932 11348 30984 11354
rect 30932 11290 30984 11296
rect 31036 11150 31064 12106
rect 31128 11694 31156 12922
rect 31220 12918 31248 13874
rect 31312 13870 31340 15558
rect 31588 15434 31616 17750
rect 32048 17746 32076 18634
rect 32036 17740 32088 17746
rect 32036 17682 32088 17688
rect 31668 17672 31720 17678
rect 31668 17614 31720 17620
rect 32034 17640 32090 17649
rect 31392 15428 31444 15434
rect 31392 15370 31444 15376
rect 31576 15428 31628 15434
rect 31576 15370 31628 15376
rect 31300 13864 31352 13870
rect 31300 13806 31352 13812
rect 31208 12912 31260 12918
rect 31208 12854 31260 12860
rect 31220 12374 31248 12854
rect 31312 12442 31340 13806
rect 31404 13258 31432 15370
rect 31392 13252 31444 13258
rect 31392 13194 31444 13200
rect 31680 12646 31708 17614
rect 32324 17610 32352 21830
rect 32876 21554 32904 22918
rect 32968 22545 32996 32710
rect 35728 32230 35756 32710
rect 35820 32230 35848 32846
rect 36280 32502 36308 32864
rect 36452 32846 36504 32852
rect 37740 32904 37792 32910
rect 37740 32846 37792 32852
rect 37556 32836 37608 32842
rect 37556 32778 37608 32784
rect 36268 32496 36320 32502
rect 36268 32438 36320 32444
rect 35716 32224 35768 32230
rect 35716 32166 35768 32172
rect 35808 32224 35860 32230
rect 35808 32166 35860 32172
rect 35728 31754 35756 32166
rect 35820 31822 35848 32166
rect 35808 31816 35860 31822
rect 35808 31758 35860 31764
rect 35716 31748 35768 31754
rect 35716 31690 35768 31696
rect 35164 31680 35216 31686
rect 35164 31622 35216 31628
rect 35176 31278 35204 31622
rect 35728 31346 35756 31690
rect 35716 31340 35768 31346
rect 35716 31282 35768 31288
rect 35164 31272 35216 31278
rect 35164 31214 35216 31220
rect 35176 30598 35204 31214
rect 35808 30728 35860 30734
rect 35808 30670 35860 30676
rect 35164 30592 35216 30598
rect 35164 30534 35216 30540
rect 35348 30592 35400 30598
rect 35348 30534 35400 30540
rect 35176 29646 35204 30534
rect 35164 29640 35216 29646
rect 35164 29582 35216 29588
rect 34796 28960 34848 28966
rect 34796 28902 34848 28908
rect 34808 28082 34836 28902
rect 35176 28422 35204 29582
rect 35360 29510 35388 30534
rect 35820 30054 35848 30670
rect 35808 30048 35860 30054
rect 35808 29990 35860 29996
rect 35820 29646 35848 29990
rect 35808 29640 35860 29646
rect 35808 29582 35860 29588
rect 35348 29504 35400 29510
rect 35348 29446 35400 29452
rect 35360 28558 35388 29446
rect 36280 29170 36308 32438
rect 37464 32224 37516 32230
rect 37464 32166 37516 32172
rect 37070 32124 37378 32133
rect 37070 32122 37076 32124
rect 37132 32122 37156 32124
rect 37212 32122 37236 32124
rect 37292 32122 37316 32124
rect 37372 32122 37378 32124
rect 37132 32070 37134 32122
rect 37314 32070 37316 32122
rect 37070 32068 37076 32070
rect 37132 32068 37156 32070
rect 37212 32068 37236 32070
rect 37292 32068 37316 32070
rect 37372 32068 37378 32070
rect 37070 32059 37378 32068
rect 37476 31822 37504 32166
rect 37568 32026 37596 32778
rect 37752 32570 37780 32846
rect 37740 32564 37792 32570
rect 37740 32506 37792 32512
rect 38568 32564 38620 32570
rect 38568 32506 38620 32512
rect 37924 32224 37976 32230
rect 37924 32166 37976 32172
rect 38476 32224 38528 32230
rect 38476 32166 38528 32172
rect 37556 32020 37608 32026
rect 37556 31962 37608 31968
rect 37464 31816 37516 31822
rect 37464 31758 37516 31764
rect 37476 31346 37504 31758
rect 37568 31482 37596 31962
rect 37936 31822 37964 32166
rect 38488 31822 38516 32166
rect 38580 32026 38608 32506
rect 38568 32020 38620 32026
rect 38568 31962 38620 31968
rect 37924 31816 37976 31822
rect 37924 31758 37976 31764
rect 38476 31816 38528 31822
rect 38476 31758 38528 31764
rect 37556 31476 37608 31482
rect 37556 31418 37608 31424
rect 37464 31340 37516 31346
rect 37464 31282 37516 31288
rect 37070 31036 37378 31045
rect 37070 31034 37076 31036
rect 37132 31034 37156 31036
rect 37212 31034 37236 31036
rect 37292 31034 37316 31036
rect 37372 31034 37378 31036
rect 37132 30982 37134 31034
rect 37314 30982 37316 31034
rect 37070 30980 37076 30982
rect 37132 30980 37156 30982
rect 37212 30980 37236 30982
rect 37292 30980 37316 30982
rect 37372 30980 37378 30982
rect 37070 30971 37378 30980
rect 37476 30734 37504 31282
rect 37568 30938 37596 31418
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 37464 30728 37516 30734
rect 37464 30670 37516 30676
rect 37372 30660 37424 30666
rect 37372 30602 37424 30608
rect 37384 30394 37412 30602
rect 37372 30388 37424 30394
rect 37372 30330 37424 30336
rect 37070 29948 37378 29957
rect 37070 29946 37076 29948
rect 37132 29946 37156 29948
rect 37212 29946 37236 29948
rect 37292 29946 37316 29948
rect 37372 29946 37378 29948
rect 37132 29894 37134 29946
rect 37314 29894 37316 29946
rect 37070 29892 37076 29894
rect 37132 29892 37156 29894
rect 37212 29892 37236 29894
rect 37292 29892 37316 29894
rect 37372 29892 37378 29894
rect 37070 29883 37378 29892
rect 37568 29850 37596 30874
rect 37936 30734 37964 31758
rect 38488 31482 38516 31758
rect 38476 31476 38528 31482
rect 38476 31418 38528 31424
rect 38488 30734 38516 31418
rect 38580 31346 38608 31962
rect 38568 31340 38620 31346
rect 38568 31282 38620 31288
rect 38580 30938 38608 31282
rect 38568 30932 38620 30938
rect 38568 30874 38620 30880
rect 37924 30728 37976 30734
rect 37924 30670 37976 30676
rect 38476 30728 38528 30734
rect 38476 30670 38528 30676
rect 37556 29844 37608 29850
rect 37556 29786 37608 29792
rect 36268 29164 36320 29170
rect 36268 29106 36320 29112
rect 36084 29028 36136 29034
rect 36084 28970 36136 28976
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 35164 28416 35216 28422
rect 35164 28358 35216 28364
rect 34796 28076 34848 28082
rect 34796 28018 34848 28024
rect 34808 27878 34836 28018
rect 35176 28014 35204 28358
rect 35360 28082 35388 28494
rect 36096 28082 36124 28970
rect 36280 28558 36308 29106
rect 37070 28860 37378 28869
rect 37070 28858 37076 28860
rect 37132 28858 37156 28860
rect 37212 28858 37236 28860
rect 37292 28858 37316 28860
rect 37372 28858 37378 28860
rect 37132 28806 37134 28858
rect 37314 28806 37316 28858
rect 37070 28804 37076 28806
rect 37132 28804 37156 28806
rect 37212 28804 37236 28806
rect 37292 28804 37316 28806
rect 37372 28804 37378 28806
rect 37070 28795 37378 28804
rect 37568 28762 37596 29786
rect 37936 29646 37964 30670
rect 38488 30394 38516 30670
rect 38476 30388 38528 30394
rect 38476 30330 38528 30336
rect 37924 29640 37976 29646
rect 37924 29582 37976 29588
rect 37556 28756 37608 28762
rect 37556 28698 37608 28704
rect 36268 28552 36320 28558
rect 36268 28494 36320 28500
rect 37568 28218 37596 28698
rect 37556 28212 37608 28218
rect 37556 28154 37608 28160
rect 35348 28076 35400 28082
rect 35348 28018 35400 28024
rect 36084 28076 36136 28082
rect 36084 28018 36136 28024
rect 35164 28008 35216 28014
rect 35164 27950 35216 27956
rect 34796 27872 34848 27878
rect 34796 27814 34848 27820
rect 34520 25220 34572 25226
rect 34520 25162 34572 25168
rect 34532 24750 34560 25162
rect 33416 24744 33468 24750
rect 33416 24686 33468 24692
rect 33600 24744 33652 24750
rect 33600 24686 33652 24692
rect 34520 24744 34572 24750
rect 34520 24686 34572 24692
rect 33428 24410 33456 24686
rect 33416 24404 33468 24410
rect 33416 24346 33468 24352
rect 33612 23769 33640 24686
rect 33968 24132 34020 24138
rect 33968 24074 34020 24080
rect 33876 23792 33928 23798
rect 33598 23760 33654 23769
rect 33876 23734 33928 23740
rect 33598 23695 33654 23704
rect 33508 22636 33560 22642
rect 33508 22578 33560 22584
rect 32954 22536 33010 22545
rect 32954 22471 33010 22480
rect 32864 21548 32916 21554
rect 32864 21490 32916 21496
rect 32404 21004 32456 21010
rect 32404 20946 32456 20952
rect 32416 20534 32444 20946
rect 32876 20806 32904 21490
rect 33416 21344 33468 21350
rect 33416 21286 33468 21292
rect 33428 20874 33456 21286
rect 33520 21146 33548 22578
rect 33888 22098 33916 23734
rect 33980 23322 34008 24074
rect 33968 23316 34020 23322
rect 33968 23258 34020 23264
rect 34060 22432 34112 22438
rect 34060 22374 34112 22380
rect 33876 22092 33928 22098
rect 34072 22094 34100 22374
rect 34072 22066 34192 22094
rect 33876 22034 33928 22040
rect 34164 22030 34192 22066
rect 34152 22024 34204 22030
rect 34152 21966 34204 21972
rect 34520 21548 34572 21554
rect 34520 21490 34572 21496
rect 33508 21140 33560 21146
rect 33508 21082 33560 21088
rect 33416 20868 33468 20874
rect 33416 20810 33468 20816
rect 32864 20800 32916 20806
rect 32864 20742 32916 20748
rect 32404 20528 32456 20534
rect 32404 20470 32456 20476
rect 32956 20528 33008 20534
rect 32956 20470 33008 20476
rect 32968 20058 32996 20470
rect 34532 20466 34560 21490
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34624 20262 34652 20878
rect 34336 20256 34388 20262
rect 34336 20198 34388 20204
rect 34612 20256 34664 20262
rect 34612 20198 34664 20204
rect 32956 20052 33008 20058
rect 32956 19994 33008 20000
rect 32496 19712 32548 19718
rect 32496 19654 32548 19660
rect 32508 19310 32536 19654
rect 32496 19304 32548 19310
rect 32496 19246 32548 19252
rect 33876 19168 33928 19174
rect 33876 19110 33928 19116
rect 33598 18728 33654 18737
rect 33598 18663 33600 18672
rect 33652 18663 33654 18672
rect 33600 18634 33652 18640
rect 33888 18358 33916 19110
rect 34348 18970 34376 20198
rect 34612 19848 34664 19854
rect 34612 19790 34664 19796
rect 34624 19378 34652 19790
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 34336 18964 34388 18970
rect 34336 18906 34388 18912
rect 33968 18760 34020 18766
rect 33968 18702 34020 18708
rect 33980 18426 34008 18702
rect 33968 18420 34020 18426
rect 33968 18362 34020 18368
rect 33876 18352 33928 18358
rect 33876 18294 33928 18300
rect 32588 18284 32640 18290
rect 32588 18226 32640 18232
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 32034 17575 32090 17584
rect 32312 17604 32364 17610
rect 31760 16516 31812 16522
rect 31760 16458 31812 16464
rect 31772 16250 31800 16458
rect 31760 16244 31812 16250
rect 31760 16186 31812 16192
rect 32048 15638 32076 17575
rect 32312 17546 32364 17552
rect 32600 17270 32628 18226
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32220 17128 32272 17134
rect 32220 17070 32272 17076
rect 32126 16144 32182 16153
rect 32126 16079 32182 16088
rect 32140 16046 32168 16079
rect 32128 16040 32180 16046
rect 32128 15982 32180 15988
rect 32036 15632 32088 15638
rect 32036 15574 32088 15580
rect 32140 15162 32168 15982
rect 32232 15638 32260 17070
rect 32600 16998 32628 17206
rect 32588 16992 32640 16998
rect 32588 16934 32640 16940
rect 33152 16794 33180 18226
rect 33980 18086 34008 18362
rect 34808 18222 34836 27814
rect 35176 27334 35204 27950
rect 36096 27674 36124 28018
rect 37070 27772 37378 27781
rect 37070 27770 37076 27772
rect 37132 27770 37156 27772
rect 37212 27770 37236 27772
rect 37292 27770 37316 27772
rect 37372 27770 37378 27772
rect 37132 27718 37134 27770
rect 37314 27718 37316 27770
rect 37070 27716 37076 27718
rect 37132 27716 37156 27718
rect 37212 27716 37236 27718
rect 37292 27716 37316 27718
rect 37372 27716 37378 27718
rect 37070 27707 37378 27716
rect 36084 27668 36136 27674
rect 36084 27610 36136 27616
rect 35164 27328 35216 27334
rect 35164 27270 35216 27276
rect 35992 25900 36044 25906
rect 35992 25842 36044 25848
rect 34980 25288 35032 25294
rect 34980 25230 35032 25236
rect 34992 24410 35020 25230
rect 36004 24818 36032 25842
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 35348 24608 35400 24614
rect 35348 24550 35400 24556
rect 34980 24404 35032 24410
rect 34980 24346 35032 24352
rect 34992 24206 35020 24346
rect 35360 24206 35388 24550
rect 36004 24410 36032 24754
rect 35992 24404 36044 24410
rect 35992 24346 36044 24352
rect 34980 24200 35032 24206
rect 34980 24142 35032 24148
rect 35348 24200 35400 24206
rect 35348 24142 35400 24148
rect 35992 23792 36044 23798
rect 35992 23734 36044 23740
rect 35900 23520 35952 23526
rect 35900 23462 35952 23468
rect 35440 23112 35492 23118
rect 35440 23054 35492 23060
rect 35072 22976 35124 22982
rect 35072 22918 35124 22924
rect 35084 22710 35112 22918
rect 35072 22704 35124 22710
rect 35072 22646 35124 22652
rect 35452 21690 35480 23054
rect 35912 22642 35940 23462
rect 36004 23322 36032 23734
rect 35992 23316 36044 23322
rect 35992 23258 36044 23264
rect 35900 22636 35952 22642
rect 35900 22578 35952 22584
rect 35912 22030 35940 22578
rect 35900 22024 35952 22030
rect 35900 21966 35952 21972
rect 35440 21684 35492 21690
rect 35440 21626 35492 21632
rect 35624 21548 35676 21554
rect 35624 21490 35676 21496
rect 35532 21072 35584 21078
rect 35532 21014 35584 21020
rect 35072 20256 35124 20262
rect 35072 20198 35124 20204
rect 35084 19242 35112 20198
rect 35348 19440 35400 19446
rect 35348 19382 35400 19388
rect 35256 19372 35308 19378
rect 35256 19314 35308 19320
rect 35072 19236 35124 19242
rect 35072 19178 35124 19184
rect 34888 18692 34940 18698
rect 34888 18634 34940 18640
rect 34900 18426 34928 18634
rect 34888 18420 34940 18426
rect 34888 18362 34940 18368
rect 35164 18352 35216 18358
rect 35164 18294 35216 18300
rect 34244 18216 34296 18222
rect 34244 18158 34296 18164
rect 34612 18216 34664 18222
rect 34612 18158 34664 18164
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34256 18086 34284 18158
rect 33232 18080 33284 18086
rect 33232 18022 33284 18028
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 34244 18080 34296 18086
rect 34244 18022 34296 18028
rect 33244 17134 33272 18022
rect 33324 17536 33376 17542
rect 33324 17478 33376 17484
rect 33232 17128 33284 17134
rect 33232 17070 33284 17076
rect 33336 16794 33364 17478
rect 33140 16788 33192 16794
rect 33140 16730 33192 16736
rect 33324 16788 33376 16794
rect 33324 16730 33376 16736
rect 33980 16658 34008 18022
rect 34060 17536 34112 17542
rect 34060 17478 34112 17484
rect 34072 16697 34100 17478
rect 34058 16688 34114 16697
rect 33968 16652 34020 16658
rect 34058 16623 34114 16632
rect 33968 16594 34020 16600
rect 33876 16448 33928 16454
rect 33876 16390 33928 16396
rect 32404 16040 32456 16046
rect 32404 15982 32456 15988
rect 33140 16040 33192 16046
rect 33140 15982 33192 15988
rect 32416 15706 32444 15982
rect 32404 15700 32456 15706
rect 32404 15642 32456 15648
rect 32220 15632 32272 15638
rect 32220 15574 32272 15580
rect 32232 15366 32260 15574
rect 33152 15502 33180 15982
rect 33888 15978 33916 16390
rect 33876 15972 33928 15978
rect 33876 15914 33928 15920
rect 33600 15564 33652 15570
rect 33600 15506 33652 15512
rect 33140 15496 33192 15502
rect 33140 15438 33192 15444
rect 32404 15428 32456 15434
rect 32404 15370 32456 15376
rect 32220 15360 32272 15366
rect 32220 15302 32272 15308
rect 32128 15156 32180 15162
rect 32128 15098 32180 15104
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32220 14816 32272 14822
rect 32220 14758 32272 14764
rect 32232 14346 32260 14758
rect 32324 14550 32352 14962
rect 32312 14544 32364 14550
rect 32312 14486 32364 14492
rect 32220 14340 32272 14346
rect 32220 14282 32272 14288
rect 32416 13802 32444 15370
rect 33612 15026 33640 15506
rect 33980 15502 34008 16594
rect 34256 16522 34284 18022
rect 34624 17542 34652 18158
rect 34704 18148 34756 18154
rect 34704 18090 34756 18096
rect 34612 17536 34664 17542
rect 34612 17478 34664 17484
rect 34716 17202 34744 18090
rect 34808 17746 34836 18158
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 34796 17264 34848 17270
rect 34796 17206 34848 17212
rect 34704 17196 34756 17202
rect 34704 17138 34756 17144
rect 34808 16590 34836 17206
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 34244 16516 34296 16522
rect 34244 16458 34296 16464
rect 34060 16448 34112 16454
rect 34060 16390 34112 16396
rect 34072 16182 34100 16390
rect 34060 16176 34112 16182
rect 34060 16118 34112 16124
rect 34888 15904 34940 15910
rect 34888 15846 34940 15852
rect 33968 15496 34020 15502
rect 33968 15438 34020 15444
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33048 14952 33100 14958
rect 33048 14894 33100 14900
rect 33232 14952 33284 14958
rect 33232 14894 33284 14900
rect 32588 14272 32640 14278
rect 32588 14214 32640 14220
rect 32600 13852 32628 14214
rect 32680 13864 32732 13870
rect 32600 13824 32680 13852
rect 32404 13796 32456 13802
rect 32404 13738 32456 13744
rect 32600 13394 32628 13824
rect 32680 13806 32732 13812
rect 32588 13388 32640 13394
rect 32588 13330 32640 13336
rect 32220 13184 32272 13190
rect 32220 13126 32272 13132
rect 32232 12782 32260 13126
rect 32220 12776 32272 12782
rect 32220 12718 32272 12724
rect 31484 12640 31536 12646
rect 31484 12582 31536 12588
rect 31668 12640 31720 12646
rect 31668 12582 31720 12588
rect 31300 12436 31352 12442
rect 31300 12378 31352 12384
rect 31392 12436 31444 12442
rect 31496 12434 31524 12582
rect 31444 12406 31524 12434
rect 31392 12378 31444 12384
rect 31208 12368 31260 12374
rect 31208 12310 31260 12316
rect 31220 12238 31248 12310
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 31404 11762 31432 12378
rect 31576 12096 31628 12102
rect 31576 12038 31628 12044
rect 31588 11762 31616 12038
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31576 11756 31628 11762
rect 31576 11698 31628 11704
rect 31668 11756 31720 11762
rect 31668 11698 31720 11704
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 31116 11688 31168 11694
rect 31116 11630 31168 11636
rect 31220 11642 31248 11698
rect 31680 11642 31708 11698
rect 31220 11614 31708 11642
rect 31668 11348 31720 11354
rect 31668 11290 31720 11296
rect 31024 11144 31076 11150
rect 31024 11086 31076 11092
rect 31680 11098 31708 11290
rect 31036 10266 31064 11086
rect 31680 11070 31800 11098
rect 31668 11008 31720 11014
rect 31668 10950 31720 10956
rect 31024 10260 31076 10266
rect 31024 10202 31076 10208
rect 31484 10260 31536 10266
rect 31484 10202 31536 10208
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 30852 9926 30880 10066
rect 30840 9920 30892 9926
rect 30840 9862 30892 9868
rect 30708 9676 30788 9704
rect 30656 9658 30708 9664
rect 30668 9518 30696 9658
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30656 9512 30708 9518
rect 30656 9454 30708 9460
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30196 6792 30248 6798
rect 30196 6734 30248 6740
rect 29736 6656 29788 6662
rect 29736 6598 29788 6604
rect 29748 6254 29776 6598
rect 29846 6556 30154 6565
rect 29846 6554 29852 6556
rect 29908 6554 29932 6556
rect 29988 6554 30012 6556
rect 30068 6554 30092 6556
rect 30148 6554 30154 6556
rect 29908 6502 29910 6554
rect 30090 6502 30092 6554
rect 29846 6500 29852 6502
rect 29908 6500 29932 6502
rect 29988 6500 30012 6502
rect 30068 6500 30092 6502
rect 30148 6500 30154 6502
rect 29846 6491 30154 6500
rect 29736 6248 29788 6254
rect 29736 6190 29788 6196
rect 30208 6118 30236 6734
rect 30196 6112 30248 6118
rect 30196 6054 30248 6060
rect 29846 5468 30154 5477
rect 29846 5466 29852 5468
rect 29908 5466 29932 5468
rect 29988 5466 30012 5468
rect 30068 5466 30092 5468
rect 30148 5466 30154 5468
rect 29908 5414 29910 5466
rect 30090 5414 30092 5466
rect 29846 5412 29852 5414
rect 29908 5412 29932 5414
rect 29988 5412 30012 5414
rect 30068 5412 30092 5414
rect 30148 5412 30154 5414
rect 29846 5403 30154 5412
rect 30300 5302 30328 8434
rect 30576 8412 30604 9454
rect 31496 8906 31524 10202
rect 31680 10198 31708 10950
rect 31772 10674 31800 11070
rect 32508 11014 32536 11698
rect 32956 11688 33008 11694
rect 32956 11630 33008 11636
rect 32588 11552 32640 11558
rect 32588 11494 32640 11500
rect 32600 11150 32628 11494
rect 32968 11354 32996 11630
rect 32956 11348 33008 11354
rect 32956 11290 33008 11296
rect 32588 11144 32640 11150
rect 32588 11086 32640 11092
rect 32496 11008 32548 11014
rect 32496 10950 32548 10956
rect 31760 10668 31812 10674
rect 31760 10610 31812 10616
rect 32588 10464 32640 10470
rect 32588 10406 32640 10412
rect 32600 10266 32628 10406
rect 32588 10260 32640 10266
rect 32588 10202 32640 10208
rect 31668 10192 31720 10198
rect 31720 10140 31892 10146
rect 31668 10134 31892 10140
rect 31680 10130 31892 10134
rect 31680 10124 31904 10130
rect 31680 10118 31852 10124
rect 31852 10066 31904 10072
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31668 9988 31720 9994
rect 31668 9930 31720 9936
rect 31680 9897 31708 9930
rect 31666 9888 31722 9897
rect 31666 9823 31722 9832
rect 31772 9450 31800 9998
rect 31944 9580 31996 9586
rect 31944 9522 31996 9528
rect 31760 9444 31812 9450
rect 31760 9386 31812 9392
rect 31576 9036 31628 9042
rect 31576 8978 31628 8984
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 30930 8528 30986 8537
rect 30840 8492 30892 8498
rect 30930 8463 30932 8472
rect 30840 8434 30892 8440
rect 30984 8463 30986 8472
rect 30932 8434 30984 8440
rect 30748 8424 30800 8430
rect 30576 8384 30748 8412
rect 30472 8356 30524 8362
rect 30472 8298 30524 8304
rect 30484 7002 30512 8298
rect 30576 7954 30604 8384
rect 30748 8366 30800 8372
rect 30852 8090 30880 8434
rect 30840 8084 30892 8090
rect 30840 8026 30892 8032
rect 30944 8022 30972 8434
rect 31114 8120 31170 8129
rect 31114 8055 31170 8064
rect 30932 8016 30984 8022
rect 30932 7958 30984 7964
rect 30564 7948 30616 7954
rect 30564 7890 30616 7896
rect 30748 7404 30800 7410
rect 30748 7346 30800 7352
rect 30562 7032 30618 7041
rect 30472 6996 30524 7002
rect 30562 6967 30618 6976
rect 30472 6938 30524 6944
rect 30576 6798 30604 6967
rect 30472 6792 30524 6798
rect 30472 6734 30524 6740
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30484 6322 30512 6734
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 30484 5234 30512 6258
rect 30668 5658 30696 6598
rect 30760 5710 30788 7346
rect 31128 7041 31156 8055
rect 31300 7812 31352 7818
rect 31300 7754 31352 7760
rect 31312 7342 31340 7754
rect 31208 7336 31260 7342
rect 31208 7278 31260 7284
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31114 7032 31170 7041
rect 31220 7002 31248 7278
rect 31114 6967 31170 6976
rect 31208 6996 31260 7002
rect 31208 6938 31260 6944
rect 30840 6792 30892 6798
rect 30840 6734 30892 6740
rect 30852 5710 30880 6734
rect 30576 5630 30696 5658
rect 30748 5704 30800 5710
rect 30748 5646 30800 5652
rect 30840 5704 30892 5710
rect 30840 5646 30892 5652
rect 31024 5704 31076 5710
rect 31024 5646 31076 5652
rect 29644 5228 29696 5234
rect 29644 5170 29696 5176
rect 30472 5228 30524 5234
rect 30472 5170 30524 5176
rect 30576 5166 30604 5630
rect 30656 5568 30708 5574
rect 30656 5510 30708 5516
rect 30668 5370 30696 5510
rect 30656 5364 30708 5370
rect 30656 5306 30708 5312
rect 31036 5234 31064 5646
rect 31024 5228 31076 5234
rect 31024 5170 31076 5176
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30564 5160 30616 5166
rect 30564 5102 30616 5108
rect 29644 4684 29696 4690
rect 29644 4626 29696 4632
rect 29184 4616 29236 4622
rect 29184 4558 29236 4564
rect 29196 3942 29224 4558
rect 29656 4486 29684 4626
rect 29644 4480 29696 4486
rect 29644 4422 29696 4428
rect 29184 3936 29236 3942
rect 29184 3878 29236 3884
rect 29196 3738 29224 3878
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 28080 3596 28132 3602
rect 28080 3538 28132 3544
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 27896 3052 27948 3058
rect 27896 2994 27948 3000
rect 29196 2990 29224 3674
rect 29656 3194 29684 4422
rect 29846 4380 30154 4389
rect 29846 4378 29852 4380
rect 29908 4378 29932 4380
rect 29988 4378 30012 4380
rect 30068 4378 30092 4380
rect 30148 4378 30154 4380
rect 29908 4326 29910 4378
rect 30090 4326 30092 4378
rect 29846 4324 29852 4326
rect 29908 4324 29932 4326
rect 29988 4324 30012 4326
rect 30068 4324 30092 4326
rect 30148 4324 30154 4326
rect 29846 4315 30154 4324
rect 30392 3670 30420 5102
rect 31404 4690 31432 8774
rect 31496 8634 31524 8842
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31588 8378 31616 8978
rect 31496 8350 31616 8378
rect 31772 8362 31800 9386
rect 31956 8974 31984 9522
rect 32770 9072 32826 9081
rect 32770 9007 32826 9016
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 32404 8968 32456 8974
rect 32404 8910 32456 8916
rect 31760 8356 31812 8362
rect 31496 5166 31524 8350
rect 31760 8298 31812 8304
rect 31576 8288 31628 8294
rect 31576 8230 31628 8236
rect 31588 7818 31616 8230
rect 31758 8120 31814 8129
rect 31758 8055 31814 8064
rect 31772 8022 31800 8055
rect 31668 8016 31720 8022
rect 31666 7984 31668 7993
rect 31760 8016 31812 8022
rect 31720 7984 31722 7993
rect 31760 7958 31812 7964
rect 31666 7919 31722 7928
rect 31576 7812 31628 7818
rect 31576 7754 31628 7760
rect 31852 7744 31904 7750
rect 31852 7686 31904 7692
rect 31576 7404 31628 7410
rect 31576 7346 31628 7352
rect 31588 7041 31616 7346
rect 31574 7032 31630 7041
rect 31864 7002 31892 7686
rect 31574 6967 31630 6976
rect 31852 6996 31904 7002
rect 31852 6938 31904 6944
rect 31574 6896 31630 6905
rect 31574 6831 31576 6840
rect 31628 6831 31630 6840
rect 31576 6802 31628 6808
rect 31484 5160 31536 5166
rect 31484 5102 31536 5108
rect 31392 4684 31444 4690
rect 31392 4626 31444 4632
rect 31496 4622 31524 5102
rect 31484 4616 31536 4622
rect 31484 4558 31536 4564
rect 31760 4548 31812 4554
rect 31760 4490 31812 4496
rect 31772 4282 31800 4490
rect 31760 4276 31812 4282
rect 31760 4218 31812 4224
rect 31956 3942 31984 8910
rect 32312 8832 32364 8838
rect 32312 8774 32364 8780
rect 32128 8560 32180 8566
rect 32128 8502 32180 8508
rect 32036 8424 32088 8430
rect 32036 8366 32088 8372
rect 32048 7886 32076 8366
rect 32036 7880 32088 7886
rect 32036 7822 32088 7828
rect 32140 7818 32168 8502
rect 32324 8498 32352 8774
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32416 8430 32444 8910
rect 32680 8900 32732 8906
rect 32680 8842 32732 8848
rect 32692 8634 32720 8842
rect 32784 8634 32812 9007
rect 33060 8634 33088 14894
rect 33140 13184 33192 13190
rect 33140 13126 33192 13132
rect 33152 12782 33180 13126
rect 33140 12776 33192 12782
rect 33140 12718 33192 12724
rect 33152 12102 33180 12718
rect 33244 12714 33272 14894
rect 33612 13938 33640 14962
rect 33980 14618 34008 15438
rect 33968 14612 34020 14618
rect 33968 14554 34020 14560
rect 33600 13932 33652 13938
rect 33600 13874 33652 13880
rect 33612 12850 33640 13874
rect 33980 13530 34008 14554
rect 34900 14006 34928 15846
rect 35176 15162 35204 18294
rect 35268 17678 35296 19314
rect 35256 17672 35308 17678
rect 35256 17614 35308 17620
rect 35268 16182 35296 17614
rect 35360 16590 35388 19382
rect 35440 19304 35492 19310
rect 35440 19246 35492 19252
rect 35452 18426 35480 19246
rect 35440 18420 35492 18426
rect 35440 18362 35492 18368
rect 35544 16590 35572 21014
rect 35636 19854 35664 21490
rect 35808 21344 35860 21350
rect 35808 21286 35860 21292
rect 35820 20534 35848 21286
rect 35808 20528 35860 20534
rect 35808 20470 35860 20476
rect 35624 19848 35676 19854
rect 35624 19790 35676 19796
rect 36096 19310 36124 27610
rect 37070 26684 37378 26693
rect 37070 26682 37076 26684
rect 37132 26682 37156 26684
rect 37212 26682 37236 26684
rect 37292 26682 37316 26684
rect 37372 26682 37378 26684
rect 37132 26630 37134 26682
rect 37314 26630 37316 26682
rect 37070 26628 37076 26630
rect 37132 26628 37156 26630
rect 37212 26628 37236 26630
rect 37292 26628 37316 26630
rect 37372 26628 37378 26630
rect 37070 26619 37378 26628
rect 37568 26314 37596 28154
rect 40960 27668 41012 27674
rect 40960 27610 41012 27616
rect 40776 26580 40828 26586
rect 40776 26522 40828 26528
rect 37648 26376 37700 26382
rect 37648 26318 37700 26324
rect 37556 26308 37608 26314
rect 37556 26250 37608 26256
rect 37070 25596 37378 25605
rect 37070 25594 37076 25596
rect 37132 25594 37156 25596
rect 37212 25594 37236 25596
rect 37292 25594 37316 25596
rect 37372 25594 37378 25596
rect 37132 25542 37134 25594
rect 37314 25542 37316 25594
rect 37070 25540 37076 25542
rect 37132 25540 37156 25542
rect 37212 25540 37236 25542
rect 37292 25540 37316 25542
rect 37372 25540 37378 25542
rect 37070 25531 37378 25540
rect 37372 24744 37424 24750
rect 37370 24712 37372 24721
rect 37424 24712 37426 24721
rect 37370 24647 37426 24656
rect 37070 24508 37378 24517
rect 37070 24506 37076 24508
rect 37132 24506 37156 24508
rect 37212 24506 37236 24508
rect 37292 24506 37316 24508
rect 37372 24506 37378 24508
rect 37132 24454 37134 24506
rect 37314 24454 37316 24506
rect 37070 24452 37076 24454
rect 37132 24452 37156 24454
rect 37212 24452 37236 24454
rect 37292 24452 37316 24454
rect 37372 24452 37378 24454
rect 37070 24443 37378 24452
rect 37556 24064 37608 24070
rect 37556 24006 37608 24012
rect 37568 23798 37596 24006
rect 37556 23792 37608 23798
rect 37556 23734 37608 23740
rect 36544 23656 36596 23662
rect 36544 23598 36596 23604
rect 36268 23180 36320 23186
rect 36268 23122 36320 23128
rect 36280 21690 36308 23122
rect 36360 23112 36412 23118
rect 36360 23054 36412 23060
rect 36268 21684 36320 21690
rect 36268 21626 36320 21632
rect 36372 21146 36400 23054
rect 36556 22574 36584 23598
rect 37070 23420 37378 23429
rect 37070 23418 37076 23420
rect 37132 23418 37156 23420
rect 37212 23418 37236 23420
rect 37292 23418 37316 23420
rect 37372 23418 37378 23420
rect 37132 23366 37134 23418
rect 37314 23366 37316 23418
rect 37070 23364 37076 23366
rect 37132 23364 37156 23366
rect 37212 23364 37236 23366
rect 37292 23364 37316 23366
rect 37372 23364 37378 23366
rect 37070 23355 37378 23364
rect 36544 22568 36596 22574
rect 36544 22510 36596 22516
rect 37070 22332 37378 22341
rect 37070 22330 37076 22332
rect 37132 22330 37156 22332
rect 37212 22330 37236 22332
rect 37292 22330 37316 22332
rect 37372 22330 37378 22332
rect 37132 22278 37134 22330
rect 37314 22278 37316 22330
rect 37070 22276 37076 22278
rect 37132 22276 37156 22278
rect 37212 22276 37236 22278
rect 37292 22276 37316 22278
rect 37372 22276 37378 22278
rect 37070 22267 37378 22276
rect 37660 22094 37688 26318
rect 39028 24812 39080 24818
rect 39028 24754 39080 24760
rect 39040 24410 39068 24754
rect 39948 24744 40000 24750
rect 39948 24686 40000 24692
rect 39120 24608 39172 24614
rect 39120 24550 39172 24556
rect 37740 24404 37792 24410
rect 37740 24346 37792 24352
rect 38568 24404 38620 24410
rect 38568 24346 38620 24352
rect 39028 24404 39080 24410
rect 39028 24346 39080 24352
rect 37752 22642 37780 24346
rect 38580 24206 38608 24346
rect 39132 24274 39160 24550
rect 39960 24410 39988 24686
rect 39948 24404 40000 24410
rect 39948 24346 40000 24352
rect 40684 24336 40736 24342
rect 40684 24278 40736 24284
rect 39120 24268 39172 24274
rect 39120 24210 39172 24216
rect 38568 24200 38620 24206
rect 38568 24142 38620 24148
rect 39132 23730 39160 24210
rect 39856 24200 39908 24206
rect 39856 24142 39908 24148
rect 38660 23724 38712 23730
rect 38660 23666 38712 23672
rect 39120 23724 39172 23730
rect 39120 23666 39172 23672
rect 38672 23322 38700 23666
rect 39868 23662 39896 24142
rect 40696 23798 40724 24278
rect 40684 23792 40736 23798
rect 40684 23734 40736 23740
rect 39856 23656 39908 23662
rect 39856 23598 39908 23604
rect 38660 23316 38712 23322
rect 38660 23258 38712 23264
rect 38384 23112 38436 23118
rect 38384 23054 38436 23060
rect 38396 22642 38424 23054
rect 40788 22710 40816 26522
rect 40776 22704 40828 22710
rect 40776 22646 40828 22652
rect 37740 22636 37792 22642
rect 37740 22578 37792 22584
rect 38384 22636 38436 22642
rect 38384 22578 38436 22584
rect 39764 22636 39816 22642
rect 39764 22578 39816 22584
rect 37752 22522 37780 22578
rect 37752 22494 37872 22522
rect 37740 22432 37792 22438
rect 37740 22374 37792 22380
rect 37568 22066 37688 22094
rect 36728 22024 36780 22030
rect 36728 21966 36780 21972
rect 36360 21140 36412 21146
rect 36360 21082 36412 21088
rect 36740 21049 36768 21966
rect 36912 21888 36964 21894
rect 36912 21830 36964 21836
rect 36820 21480 36872 21486
rect 36820 21422 36872 21428
rect 36726 21040 36782 21049
rect 36726 20975 36782 20984
rect 36544 20936 36596 20942
rect 36544 20878 36596 20884
rect 36556 20806 36584 20878
rect 36544 20800 36596 20806
rect 36544 20742 36596 20748
rect 36268 19712 36320 19718
rect 36268 19654 36320 19660
rect 36280 19514 36308 19654
rect 36268 19508 36320 19514
rect 36268 19450 36320 19456
rect 36084 19304 36136 19310
rect 36084 19246 36136 19252
rect 36096 18766 36124 19246
rect 36084 18760 36136 18766
rect 36084 18702 36136 18708
rect 36280 18698 36308 19450
rect 36268 18692 36320 18698
rect 36268 18634 36320 18640
rect 36544 18352 36596 18358
rect 36544 18294 36596 18300
rect 36452 18216 36504 18222
rect 36452 18158 36504 18164
rect 36268 17740 36320 17746
rect 36268 17682 36320 17688
rect 35900 17672 35952 17678
rect 35900 17614 35952 17620
rect 35808 17604 35860 17610
rect 35808 17546 35860 17552
rect 35820 17270 35848 17546
rect 35808 17264 35860 17270
rect 35808 17206 35860 17212
rect 35912 16794 35940 17614
rect 36176 17604 36228 17610
rect 36176 17546 36228 17552
rect 35992 17128 36044 17134
rect 35992 17070 36044 17076
rect 35900 16788 35952 16794
rect 35900 16730 35952 16736
rect 35808 16720 35860 16726
rect 35808 16662 35860 16668
rect 35348 16584 35400 16590
rect 35348 16526 35400 16532
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 35256 16176 35308 16182
rect 35256 16118 35308 16124
rect 35268 15434 35296 16118
rect 35820 16046 35848 16662
rect 35808 16040 35860 16046
rect 35808 15982 35860 15988
rect 35256 15428 35308 15434
rect 35256 15370 35308 15376
rect 35164 15156 35216 15162
rect 35164 15098 35216 15104
rect 35268 15094 35296 15370
rect 36004 15162 36032 17070
rect 36084 16992 36136 16998
rect 36084 16934 36136 16940
rect 36096 15638 36124 16934
rect 36188 16046 36216 17546
rect 36280 16114 36308 17682
rect 36464 17202 36492 18158
rect 36452 17196 36504 17202
rect 36452 17138 36504 17144
rect 36360 17060 36412 17066
rect 36360 17002 36412 17008
rect 36372 16658 36400 17002
rect 36360 16652 36412 16658
rect 36360 16594 36412 16600
rect 36268 16108 36320 16114
rect 36268 16050 36320 16056
rect 36176 16040 36228 16046
rect 36176 15982 36228 15988
rect 36360 15700 36412 15706
rect 36360 15642 36412 15648
rect 36084 15632 36136 15638
rect 36084 15574 36136 15580
rect 35440 15156 35492 15162
rect 35440 15098 35492 15104
rect 35992 15156 36044 15162
rect 35992 15098 36044 15104
rect 35256 15088 35308 15094
rect 35256 15030 35308 15036
rect 34244 14000 34296 14006
rect 34244 13942 34296 13948
rect 34888 14000 34940 14006
rect 34888 13942 34940 13948
rect 34256 13870 34284 13942
rect 34244 13864 34296 13870
rect 34900 13852 34928 13942
rect 34244 13806 34296 13812
rect 34808 13824 34928 13852
rect 33968 13524 34020 13530
rect 33968 13466 34020 13472
rect 33692 13252 33744 13258
rect 33692 13194 33744 13200
rect 33600 12844 33652 12850
rect 33600 12786 33652 12792
rect 33232 12708 33284 12714
rect 33232 12650 33284 12656
rect 33704 12442 33732 13194
rect 34808 13190 34836 13824
rect 34796 13184 34848 13190
rect 34796 13126 34848 13132
rect 34808 12918 34836 13126
rect 35348 12980 35400 12986
rect 35452 12968 35480 15098
rect 36268 13320 36320 13326
rect 36268 13262 36320 13268
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 35544 12986 35572 13194
rect 35400 12940 35480 12968
rect 35348 12922 35400 12928
rect 34796 12912 34848 12918
rect 34796 12854 34848 12860
rect 33784 12844 33836 12850
rect 33784 12786 33836 12792
rect 33692 12436 33744 12442
rect 33692 12378 33744 12384
rect 33416 12300 33468 12306
rect 33416 12242 33468 12248
rect 33140 12096 33192 12102
rect 33140 12038 33192 12044
rect 33152 9994 33180 12038
rect 33428 11898 33456 12242
rect 33704 12238 33732 12378
rect 33692 12232 33744 12238
rect 33692 12174 33744 12180
rect 33416 11892 33468 11898
rect 33416 11834 33468 11840
rect 33600 11756 33652 11762
rect 33600 11698 33652 11704
rect 33612 11082 33640 11698
rect 33600 11076 33652 11082
rect 33600 11018 33652 11024
rect 33796 10742 33824 12786
rect 34060 12776 34112 12782
rect 34060 12718 34112 12724
rect 34072 12374 34100 12718
rect 35452 12646 35480 12940
rect 35532 12980 35584 12986
rect 35532 12922 35584 12928
rect 35544 12782 35572 12922
rect 35992 12844 36044 12850
rect 35992 12786 36044 12792
rect 35532 12776 35584 12782
rect 35532 12718 35584 12724
rect 35440 12640 35492 12646
rect 35440 12582 35492 12588
rect 34060 12368 34112 12374
rect 34060 12310 34112 12316
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 34520 12164 34572 12170
rect 34520 12106 34572 12112
rect 34532 11762 34560 12106
rect 34808 11898 34836 12242
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 34900 11762 34928 12174
rect 35452 11762 35480 12582
rect 35544 11898 35572 12718
rect 35900 12300 35952 12306
rect 35900 12242 35952 12248
rect 35532 11892 35584 11898
rect 35532 11834 35584 11840
rect 35912 11762 35940 12242
rect 36004 11830 36032 12786
rect 36280 12238 36308 13262
rect 36372 12306 36400 15642
rect 36464 15026 36492 17138
rect 36556 15706 36584 18294
rect 36832 17882 36860 21422
rect 36924 18902 36952 21830
rect 37004 21548 37056 21554
rect 37004 21490 37056 21496
rect 37016 21298 37044 21490
rect 37004 21270 37044 21298
rect 37004 21162 37032 21270
rect 37070 21244 37378 21253
rect 37070 21242 37076 21244
rect 37132 21242 37156 21244
rect 37212 21242 37236 21244
rect 37292 21242 37316 21244
rect 37372 21242 37378 21244
rect 37132 21190 37134 21242
rect 37314 21190 37316 21242
rect 37070 21188 37076 21190
rect 37132 21188 37156 21190
rect 37212 21188 37236 21190
rect 37292 21188 37316 21190
rect 37372 21188 37378 21190
rect 37070 21179 37378 21188
rect 37004 21134 37044 21162
rect 37016 20942 37044 21134
rect 37004 20936 37056 20942
rect 37004 20878 37056 20884
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37070 20156 37378 20165
rect 37070 20154 37076 20156
rect 37132 20154 37156 20156
rect 37212 20154 37236 20156
rect 37292 20154 37316 20156
rect 37372 20154 37378 20156
rect 37132 20102 37134 20154
rect 37314 20102 37316 20154
rect 37070 20100 37076 20102
rect 37132 20100 37156 20102
rect 37212 20100 37236 20102
rect 37292 20100 37316 20102
rect 37372 20100 37378 20102
rect 37070 20091 37378 20100
rect 37476 19378 37504 20402
rect 37464 19372 37516 19378
rect 37464 19314 37516 19320
rect 37070 19068 37378 19077
rect 37070 19066 37076 19068
rect 37132 19066 37156 19068
rect 37212 19066 37236 19068
rect 37292 19066 37316 19068
rect 37372 19066 37378 19068
rect 37132 19014 37134 19066
rect 37314 19014 37316 19066
rect 37070 19012 37076 19014
rect 37132 19012 37156 19014
rect 37212 19012 37236 19014
rect 37292 19012 37316 19014
rect 37372 19012 37378 19014
rect 37070 19003 37378 19012
rect 36912 18896 36964 18902
rect 36912 18838 36964 18844
rect 37070 17980 37378 17989
rect 37070 17978 37076 17980
rect 37132 17978 37156 17980
rect 37212 17978 37236 17980
rect 37292 17978 37316 17980
rect 37372 17978 37378 17980
rect 37132 17926 37134 17978
rect 37314 17926 37316 17978
rect 37070 17924 37076 17926
rect 37132 17924 37156 17926
rect 37212 17924 37236 17926
rect 37292 17924 37316 17926
rect 37372 17924 37378 17926
rect 37070 17915 37378 17924
rect 36820 17876 36872 17882
rect 36820 17818 36872 17824
rect 37188 17808 37240 17814
rect 37188 17750 37240 17756
rect 37200 17338 37228 17750
rect 37188 17332 37240 17338
rect 37188 17274 37240 17280
rect 37070 16892 37378 16901
rect 37070 16890 37076 16892
rect 37132 16890 37156 16892
rect 37212 16890 37236 16892
rect 37292 16890 37316 16892
rect 37372 16890 37378 16892
rect 37132 16838 37134 16890
rect 37314 16838 37316 16890
rect 37070 16836 37076 16838
rect 37132 16836 37156 16838
rect 37212 16836 37236 16838
rect 37292 16836 37316 16838
rect 37372 16836 37378 16838
rect 37070 16827 37378 16836
rect 37070 15804 37378 15813
rect 37070 15802 37076 15804
rect 37132 15802 37156 15804
rect 37212 15802 37236 15804
rect 37292 15802 37316 15804
rect 37372 15802 37378 15804
rect 37132 15750 37134 15802
rect 37314 15750 37316 15802
rect 37070 15748 37076 15750
rect 37132 15748 37156 15750
rect 37212 15748 37236 15750
rect 37292 15748 37316 15750
rect 37372 15748 37378 15750
rect 37070 15739 37378 15748
rect 36544 15700 36596 15706
rect 36544 15642 36596 15648
rect 36544 15360 36596 15366
rect 36544 15302 36596 15308
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 36556 14346 36584 15302
rect 36636 14816 36688 14822
rect 36636 14758 36688 14764
rect 36648 14482 36676 14758
rect 37070 14716 37378 14725
rect 37070 14714 37076 14716
rect 37132 14714 37156 14716
rect 37212 14714 37236 14716
rect 37292 14714 37316 14716
rect 37372 14714 37378 14716
rect 37132 14662 37134 14714
rect 37314 14662 37316 14714
rect 37070 14660 37076 14662
rect 37132 14660 37156 14662
rect 37212 14660 37236 14662
rect 37292 14660 37316 14662
rect 37372 14660 37378 14662
rect 37070 14651 37378 14660
rect 37096 14612 37148 14618
rect 37096 14554 37148 14560
rect 36636 14476 36688 14482
rect 36636 14418 36688 14424
rect 36544 14340 36596 14346
rect 36544 14282 36596 14288
rect 37108 14278 37136 14554
rect 37096 14272 37148 14278
rect 37096 14214 37148 14220
rect 37070 13628 37378 13637
rect 37070 13626 37076 13628
rect 37132 13626 37156 13628
rect 37212 13626 37236 13628
rect 37292 13626 37316 13628
rect 37372 13626 37378 13628
rect 37132 13574 37134 13626
rect 37314 13574 37316 13626
rect 37070 13572 37076 13574
rect 37132 13572 37156 13574
rect 37212 13572 37236 13574
rect 37292 13572 37316 13574
rect 37372 13572 37378 13574
rect 37070 13563 37378 13572
rect 36912 13388 36964 13394
rect 36912 13330 36964 13336
rect 36924 12374 36952 13330
rect 37464 12776 37516 12782
rect 37464 12718 37516 12724
rect 37070 12540 37378 12549
rect 37070 12538 37076 12540
rect 37132 12538 37156 12540
rect 37212 12538 37236 12540
rect 37292 12538 37316 12540
rect 37372 12538 37378 12540
rect 37132 12486 37134 12538
rect 37314 12486 37316 12538
rect 37070 12484 37076 12486
rect 37132 12484 37156 12486
rect 37212 12484 37236 12486
rect 37292 12484 37316 12486
rect 37372 12484 37378 12486
rect 37070 12475 37378 12484
rect 36912 12368 36964 12374
rect 36912 12310 36964 12316
rect 36360 12300 36412 12306
rect 36360 12242 36412 12248
rect 36268 12232 36320 12238
rect 36268 12174 36320 12180
rect 35992 11824 36044 11830
rect 35992 11766 36044 11772
rect 34520 11756 34572 11762
rect 34520 11698 34572 11704
rect 34888 11756 34940 11762
rect 34888 11698 34940 11704
rect 35440 11756 35492 11762
rect 35440 11698 35492 11704
rect 35900 11756 35952 11762
rect 35900 11698 35952 11704
rect 34532 11354 34560 11698
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 36268 11552 36320 11558
rect 36268 11494 36320 11500
rect 34520 11348 34572 11354
rect 34520 11290 34572 11296
rect 35360 11218 35388 11494
rect 35348 11212 35400 11218
rect 35348 11154 35400 11160
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 35072 11144 35124 11150
rect 35072 11086 35124 11092
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 33796 10282 33824 10678
rect 33704 10254 33824 10282
rect 33324 10192 33376 10198
rect 33324 10134 33376 10140
rect 33140 9988 33192 9994
rect 33140 9930 33192 9936
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 32404 8424 32456 8430
rect 32404 8366 32456 8372
rect 32232 8090 32260 8366
rect 32220 8084 32272 8090
rect 32220 8026 32272 8032
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32128 7812 32180 7818
rect 32128 7754 32180 7760
rect 32232 6866 32260 7890
rect 32220 6860 32272 6866
rect 32220 6802 32272 6808
rect 32416 6254 32444 8366
rect 33048 8084 33100 8090
rect 33048 8026 33100 8032
rect 33060 7954 33088 8026
rect 33048 7948 33100 7954
rect 33048 7890 33100 7896
rect 32496 7880 32548 7886
rect 32496 7822 32548 7828
rect 32404 6248 32456 6254
rect 32404 6190 32456 6196
rect 32220 6112 32272 6118
rect 32220 6054 32272 6060
rect 32232 5642 32260 6054
rect 32312 5908 32364 5914
rect 32312 5850 32364 5856
rect 32324 5710 32352 5850
rect 32416 5778 32444 6190
rect 32508 5914 32536 7822
rect 32680 7812 32732 7818
rect 32680 7754 32732 7760
rect 32692 7546 32720 7754
rect 32680 7540 32732 7546
rect 32680 7482 32732 7488
rect 33046 7440 33102 7449
rect 33046 7375 33048 7384
rect 33100 7375 33102 7384
rect 33048 7346 33100 7352
rect 32588 6112 32640 6118
rect 32588 6054 32640 6060
rect 32496 5908 32548 5914
rect 32496 5850 32548 5856
rect 32404 5772 32456 5778
rect 32404 5714 32456 5720
rect 32312 5704 32364 5710
rect 32312 5646 32364 5652
rect 32220 5636 32272 5642
rect 32220 5578 32272 5584
rect 32324 5234 32352 5646
rect 32312 5228 32364 5234
rect 32312 5170 32364 5176
rect 32036 5160 32088 5166
rect 32036 5102 32088 5108
rect 32048 4622 32076 5102
rect 32128 5024 32180 5030
rect 32128 4966 32180 4972
rect 32036 4616 32088 4622
rect 32036 4558 32088 4564
rect 32140 4146 32168 4966
rect 32416 4146 32444 5714
rect 32600 5234 32628 6054
rect 32772 5772 32824 5778
rect 32772 5714 32824 5720
rect 32784 5642 32812 5714
rect 32772 5636 32824 5642
rect 32772 5578 32824 5584
rect 32496 5228 32548 5234
rect 32496 5170 32548 5176
rect 32588 5228 32640 5234
rect 32588 5170 32640 5176
rect 32508 4826 32536 5170
rect 33048 5092 33100 5098
rect 33048 5034 33100 5040
rect 32496 4820 32548 4826
rect 32496 4762 32548 4768
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 32404 4140 32456 4146
rect 32404 4082 32456 4088
rect 31944 3936 31996 3942
rect 31944 3878 31996 3884
rect 30380 3664 30432 3670
rect 30380 3606 30432 3612
rect 29846 3292 30154 3301
rect 29846 3290 29852 3292
rect 29908 3290 29932 3292
rect 29988 3290 30012 3292
rect 30068 3290 30092 3292
rect 30148 3290 30154 3292
rect 29908 3238 29910 3290
rect 30090 3238 30092 3290
rect 29846 3236 29852 3238
rect 29908 3236 29932 3238
rect 29988 3236 30012 3238
rect 30068 3236 30092 3238
rect 30148 3236 30154 3238
rect 29846 3227 30154 3236
rect 29644 3188 29696 3194
rect 29644 3130 29696 3136
rect 32416 3058 32444 4082
rect 32588 3936 32640 3942
rect 32588 3878 32640 3884
rect 32600 3738 32628 3878
rect 32588 3732 32640 3738
rect 32588 3674 32640 3680
rect 33060 3398 33088 5034
rect 33152 4826 33180 9930
rect 33336 9382 33364 10134
rect 33704 10130 33732 10254
rect 35084 10130 35112 11086
rect 35452 11082 35480 11154
rect 35440 11076 35492 11082
rect 35440 11018 35492 11024
rect 33692 10124 33744 10130
rect 33692 10066 33744 10072
rect 34704 10124 34756 10130
rect 34704 10066 34756 10072
rect 35072 10124 35124 10130
rect 35072 10066 35124 10072
rect 33704 9586 33732 10066
rect 34612 9988 34664 9994
rect 34612 9930 34664 9936
rect 34336 9920 34388 9926
rect 34336 9862 34388 9868
rect 33692 9580 33744 9586
rect 33692 9522 33744 9528
rect 33968 9512 34020 9518
rect 33968 9454 34020 9460
rect 33692 9444 33744 9450
rect 33692 9386 33744 9392
rect 33324 9376 33376 9382
rect 33324 9318 33376 9324
rect 33704 9110 33732 9386
rect 33980 9178 34008 9454
rect 33968 9172 34020 9178
rect 33968 9114 34020 9120
rect 34152 9172 34204 9178
rect 34152 9114 34204 9120
rect 33692 9104 33744 9110
rect 33692 9046 33744 9052
rect 34164 8294 34192 9114
rect 34348 8906 34376 9862
rect 34624 9722 34652 9930
rect 34612 9716 34664 9722
rect 34612 9658 34664 9664
rect 34336 8900 34388 8906
rect 34336 8842 34388 8848
rect 34428 8900 34480 8906
rect 34428 8842 34480 8848
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 34152 8288 34204 8294
rect 34152 8230 34204 8236
rect 34256 7954 34284 8774
rect 34348 8634 34376 8842
rect 34336 8628 34388 8634
rect 34336 8570 34388 8576
rect 34244 7948 34296 7954
rect 34244 7890 34296 7896
rect 33692 7880 33744 7886
rect 33690 7848 33692 7857
rect 33744 7848 33746 7857
rect 33690 7783 33746 7792
rect 33784 7744 33836 7750
rect 33784 7686 33836 7692
rect 34336 7744 34388 7750
rect 34336 7686 34388 7692
rect 33600 7268 33652 7274
rect 33600 7210 33652 7216
rect 33612 6390 33640 7210
rect 33796 7002 33824 7686
rect 34244 7404 34296 7410
rect 34244 7346 34296 7352
rect 33784 6996 33836 7002
rect 33784 6938 33836 6944
rect 34256 6866 34284 7346
rect 34348 7342 34376 7686
rect 34440 7546 34468 8842
rect 34520 8288 34572 8294
rect 34520 8230 34572 8236
rect 34532 7886 34560 8230
rect 34716 7954 34744 10066
rect 36280 9994 36308 11494
rect 37070 11452 37378 11461
rect 37070 11450 37076 11452
rect 37132 11450 37156 11452
rect 37212 11450 37236 11452
rect 37292 11450 37316 11452
rect 37372 11450 37378 11452
rect 37132 11398 37134 11450
rect 37314 11398 37316 11450
rect 37070 11396 37076 11398
rect 37132 11396 37156 11398
rect 37212 11396 37236 11398
rect 37292 11396 37316 11398
rect 37372 11396 37378 11398
rect 37070 11387 37378 11396
rect 36912 11212 36964 11218
rect 36912 11154 36964 11160
rect 36636 11076 36688 11082
rect 36636 11018 36688 11024
rect 36648 10810 36676 11018
rect 36636 10804 36688 10810
rect 36636 10746 36688 10752
rect 36924 10169 36952 11154
rect 37280 11076 37332 11082
rect 37280 11018 37332 11024
rect 37292 10674 37320 11018
rect 37280 10668 37332 10674
rect 37280 10610 37332 10616
rect 37476 10538 37504 12718
rect 37568 11336 37596 22066
rect 37752 21962 37780 22374
rect 37740 21956 37792 21962
rect 37740 21898 37792 21904
rect 37844 21146 37872 22494
rect 38752 22432 38804 22438
rect 38752 22374 38804 22380
rect 39212 22432 39264 22438
rect 39212 22374 39264 22380
rect 38568 21888 38620 21894
rect 38568 21830 38620 21836
rect 38580 21622 38608 21830
rect 38568 21616 38620 21622
rect 38568 21558 38620 21564
rect 38016 21548 38068 21554
rect 38016 21490 38068 21496
rect 38028 21457 38056 21490
rect 38014 21448 38070 21457
rect 38014 21383 38070 21392
rect 37832 21140 37884 21146
rect 37832 21082 37884 21088
rect 37924 20936 37976 20942
rect 37924 20878 37976 20884
rect 37936 20806 37964 20878
rect 37924 20800 37976 20806
rect 37924 20742 37976 20748
rect 38028 19854 38056 21383
rect 38476 20800 38528 20806
rect 38476 20742 38528 20748
rect 38488 19854 38516 20742
rect 38764 20534 38792 22374
rect 39224 22234 39252 22374
rect 39212 22228 39264 22234
rect 39212 22170 39264 22176
rect 39304 22024 39356 22030
rect 39304 21966 39356 21972
rect 39316 21486 39344 21966
rect 39488 21888 39540 21894
rect 39488 21830 39540 21836
rect 39304 21480 39356 21486
rect 39304 21422 39356 21428
rect 38752 20528 38804 20534
rect 38752 20470 38804 20476
rect 39500 20398 39528 21830
rect 39776 21690 39804 22578
rect 40788 22166 40816 22646
rect 40972 22642 41000 27610
rect 42708 23656 42760 23662
rect 42708 23598 42760 23604
rect 42720 23186 42748 23598
rect 42524 23180 42576 23186
rect 42524 23122 42576 23128
rect 42708 23180 42760 23186
rect 42708 23122 42760 23128
rect 42536 22642 42564 23122
rect 43352 23112 43404 23118
rect 43352 23054 43404 23060
rect 43364 22642 43392 23054
rect 40960 22636 41012 22642
rect 40960 22578 41012 22584
rect 42524 22636 42576 22642
rect 42524 22578 42576 22584
rect 43352 22636 43404 22642
rect 43352 22578 43404 22584
rect 41880 22568 41932 22574
rect 41880 22510 41932 22516
rect 40776 22160 40828 22166
rect 40776 22102 40828 22108
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 39764 21684 39816 21690
rect 39764 21626 39816 21632
rect 40052 20942 40080 21966
rect 40408 21548 40460 21554
rect 40460 21508 40632 21536
rect 40408 21490 40460 21496
rect 40604 21078 40632 21508
rect 40592 21072 40644 21078
rect 40592 21014 40644 21020
rect 39948 20936 40000 20942
rect 39948 20878 40000 20884
rect 40040 20936 40092 20942
rect 40040 20878 40092 20884
rect 39960 20602 39988 20878
rect 39948 20596 40000 20602
rect 39948 20538 40000 20544
rect 39488 20392 39540 20398
rect 39488 20334 39540 20340
rect 39396 20256 39448 20262
rect 39396 20198 39448 20204
rect 38844 20052 38896 20058
rect 38844 19994 38896 20000
rect 38016 19848 38068 19854
rect 38016 19790 38068 19796
rect 38476 19848 38528 19854
rect 38476 19790 38528 19796
rect 38384 19304 38436 19310
rect 38384 19246 38436 19252
rect 38396 18358 38424 19246
rect 38384 18352 38436 18358
rect 38384 18294 38436 18300
rect 38488 18290 38516 19790
rect 38752 19780 38804 19786
rect 38752 19722 38804 19728
rect 38764 18970 38792 19722
rect 38856 19718 38884 19994
rect 39210 19816 39266 19825
rect 39408 19786 39436 20198
rect 40052 20058 40080 20878
rect 40604 20466 40632 21014
rect 41328 20800 41380 20806
rect 41328 20742 41380 20748
rect 40316 20460 40368 20466
rect 40316 20402 40368 20408
rect 40592 20460 40644 20466
rect 40592 20402 40644 20408
rect 40132 20256 40184 20262
rect 40132 20198 40184 20204
rect 40040 20052 40092 20058
rect 40040 19994 40092 20000
rect 39210 19751 39212 19760
rect 39264 19751 39266 19760
rect 39396 19780 39448 19786
rect 39212 19722 39264 19728
rect 39396 19722 39448 19728
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 39224 19378 39252 19722
rect 39212 19372 39264 19378
rect 39212 19314 39264 19320
rect 38752 18964 38804 18970
rect 38752 18906 38804 18912
rect 38476 18284 38528 18290
rect 38476 18226 38528 18232
rect 38108 18216 38160 18222
rect 38108 18158 38160 18164
rect 38842 18184 38898 18193
rect 38120 17678 38148 18158
rect 38842 18119 38898 18128
rect 38292 17876 38344 17882
rect 38292 17818 38344 17824
rect 38108 17672 38160 17678
rect 38106 17640 38108 17649
rect 38160 17640 38162 17649
rect 38106 17575 38162 17584
rect 38304 17542 38332 17818
rect 38856 17610 38884 18119
rect 38936 17740 38988 17746
rect 38936 17682 38988 17688
rect 38844 17604 38896 17610
rect 38844 17546 38896 17552
rect 38292 17536 38344 17542
rect 38292 17478 38344 17484
rect 38568 17332 38620 17338
rect 38568 17274 38620 17280
rect 38580 17218 38608 17274
rect 38856 17270 38884 17546
rect 38844 17264 38896 17270
rect 38658 17232 38714 17241
rect 38580 17190 38658 17218
rect 38844 17206 38896 17212
rect 38658 17167 38714 17176
rect 38568 17128 38620 17134
rect 38568 17070 38620 17076
rect 38292 16992 38344 16998
rect 38292 16934 38344 16940
rect 38304 16658 38332 16934
rect 37648 16652 37700 16658
rect 37648 16594 37700 16600
rect 38292 16652 38344 16658
rect 38292 16594 38344 16600
rect 37660 16250 37688 16594
rect 37648 16244 37700 16250
rect 37648 16186 37700 16192
rect 38580 16114 38608 17070
rect 38568 16108 38620 16114
rect 38568 16050 38620 16056
rect 38844 15972 38896 15978
rect 38844 15914 38896 15920
rect 38568 15904 38620 15910
rect 38568 15846 38620 15852
rect 38580 15745 38608 15846
rect 38566 15736 38622 15745
rect 38566 15671 38622 15680
rect 38856 15570 38884 15914
rect 38660 15564 38712 15570
rect 38660 15506 38712 15512
rect 38844 15564 38896 15570
rect 38844 15506 38896 15512
rect 37648 15496 37700 15502
rect 37648 15438 37700 15444
rect 37660 14414 37688 15438
rect 38384 15428 38436 15434
rect 38384 15370 38436 15376
rect 38292 14816 38344 14822
rect 38292 14758 38344 14764
rect 38304 14414 38332 14758
rect 37648 14408 37700 14414
rect 37648 14350 37700 14356
rect 38292 14408 38344 14414
rect 38292 14350 38344 14356
rect 38200 13184 38252 13190
rect 38200 13126 38252 13132
rect 37648 12708 37700 12714
rect 37648 12650 37700 12656
rect 37660 11694 37688 12650
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 38120 11898 38148 12174
rect 38108 11892 38160 11898
rect 38108 11834 38160 11840
rect 37832 11824 37884 11830
rect 37884 11784 37964 11812
rect 37832 11766 37884 11772
rect 37648 11688 37700 11694
rect 37648 11630 37700 11636
rect 37568 11308 37872 11336
rect 37738 10704 37794 10713
rect 37738 10639 37740 10648
rect 37792 10639 37794 10648
rect 37740 10610 37792 10616
rect 37464 10532 37516 10538
rect 37464 10474 37516 10480
rect 37070 10364 37378 10373
rect 37070 10362 37076 10364
rect 37132 10362 37156 10364
rect 37212 10362 37236 10364
rect 37292 10362 37316 10364
rect 37372 10362 37378 10364
rect 37132 10310 37134 10362
rect 37314 10310 37316 10362
rect 37070 10308 37076 10310
rect 37132 10308 37156 10310
rect 37212 10308 37236 10310
rect 37292 10308 37316 10310
rect 37372 10308 37378 10310
rect 37070 10299 37378 10308
rect 36910 10160 36966 10169
rect 36910 10095 36912 10104
rect 36964 10095 36966 10104
rect 36912 10066 36964 10072
rect 36268 9988 36320 9994
rect 36268 9930 36320 9936
rect 36280 9722 36308 9930
rect 36268 9716 36320 9722
rect 36268 9658 36320 9664
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 36912 9580 36964 9586
rect 36912 9522 36964 9528
rect 35072 9444 35124 9450
rect 35072 9386 35124 9392
rect 35900 9444 35952 9450
rect 35900 9386 35952 9392
rect 35084 9110 35112 9386
rect 35072 9104 35124 9110
rect 35072 9046 35124 9052
rect 34888 9036 34940 9042
rect 34888 8978 34940 8984
rect 34900 8430 34928 8978
rect 35440 8900 35492 8906
rect 35440 8842 35492 8848
rect 35072 8832 35124 8838
rect 35072 8774 35124 8780
rect 34888 8424 34940 8430
rect 34888 8366 34940 8372
rect 34704 7948 34756 7954
rect 34704 7890 34756 7896
rect 34520 7880 34572 7886
rect 34520 7822 34572 7828
rect 34428 7540 34480 7546
rect 34428 7482 34480 7488
rect 34336 7336 34388 7342
rect 34336 7278 34388 7284
rect 34244 6860 34296 6866
rect 34244 6802 34296 6808
rect 34440 6798 34468 7482
rect 34532 6798 34560 7822
rect 34704 7200 34756 7206
rect 34704 7142 34756 7148
rect 34716 7002 34744 7142
rect 34704 6996 34756 7002
rect 34704 6938 34756 6944
rect 35084 6934 35112 8774
rect 35452 8566 35480 8842
rect 35440 8560 35492 8566
rect 35440 8502 35492 8508
rect 35072 6928 35124 6934
rect 35072 6870 35124 6876
rect 34428 6792 34480 6798
rect 34428 6734 34480 6740
rect 34520 6792 34572 6798
rect 34520 6734 34572 6740
rect 35072 6792 35124 6798
rect 35072 6734 35124 6740
rect 34440 6458 34468 6734
rect 34428 6452 34480 6458
rect 34428 6394 34480 6400
rect 33600 6384 33652 6390
rect 33600 6326 33652 6332
rect 33232 6316 33284 6322
rect 33284 6276 33364 6304
rect 33232 6258 33284 6264
rect 33232 6180 33284 6186
rect 33232 6122 33284 6128
rect 33244 5166 33272 6122
rect 33336 5370 33364 6276
rect 35084 5846 35112 6734
rect 35912 6390 35940 9386
rect 36004 8634 36032 9522
rect 36924 8838 36952 9522
rect 37070 9276 37378 9285
rect 37070 9274 37076 9276
rect 37132 9274 37156 9276
rect 37212 9274 37236 9276
rect 37292 9274 37316 9276
rect 37372 9274 37378 9276
rect 37132 9222 37134 9274
rect 37314 9222 37316 9274
rect 37070 9220 37076 9222
rect 37132 9220 37156 9222
rect 37212 9220 37236 9222
rect 37292 9220 37316 9222
rect 37372 9220 37378 9222
rect 37070 9211 37378 9220
rect 36912 8832 36964 8838
rect 36912 8774 36964 8780
rect 37740 8832 37792 8838
rect 37740 8774 37792 8780
rect 35992 8628 36044 8634
rect 35992 8570 36044 8576
rect 36004 7818 36032 8570
rect 36924 8498 36952 8774
rect 36912 8492 36964 8498
rect 36912 8434 36964 8440
rect 36924 8090 36952 8434
rect 37464 8288 37516 8294
rect 37464 8230 37516 8236
rect 37070 8188 37378 8197
rect 37070 8186 37076 8188
rect 37132 8186 37156 8188
rect 37212 8186 37236 8188
rect 37292 8186 37316 8188
rect 37372 8186 37378 8188
rect 37132 8134 37134 8186
rect 37314 8134 37316 8186
rect 37070 8132 37076 8134
rect 37132 8132 37156 8134
rect 37212 8132 37236 8134
rect 37292 8132 37316 8134
rect 37372 8132 37378 8134
rect 37070 8123 37378 8132
rect 36912 8084 36964 8090
rect 36912 8026 36964 8032
rect 37476 8022 37504 8230
rect 37464 8016 37516 8022
rect 37464 7958 37516 7964
rect 35992 7812 36044 7818
rect 35992 7754 36044 7760
rect 37752 7410 37780 8774
rect 37740 7404 37792 7410
rect 37740 7346 37792 7352
rect 36728 7268 36780 7274
rect 36728 7210 36780 7216
rect 36740 6458 36768 7210
rect 37070 7100 37378 7109
rect 37070 7098 37076 7100
rect 37132 7098 37156 7100
rect 37212 7098 37236 7100
rect 37292 7098 37316 7100
rect 37372 7098 37378 7100
rect 37132 7046 37134 7098
rect 37314 7046 37316 7098
rect 37070 7044 37076 7046
rect 37132 7044 37156 7046
rect 37212 7044 37236 7046
rect 37292 7044 37316 7046
rect 37372 7044 37378 7046
rect 37070 7035 37378 7044
rect 36728 6452 36780 6458
rect 36728 6394 36780 6400
rect 35900 6384 35952 6390
rect 35900 6326 35952 6332
rect 35072 5840 35124 5846
rect 35072 5782 35124 5788
rect 34336 5636 34388 5642
rect 34336 5578 34388 5584
rect 33324 5364 33376 5370
rect 33324 5306 33376 5312
rect 34348 5302 34376 5578
rect 34336 5296 34388 5302
rect 34336 5238 34388 5244
rect 35084 5166 35112 5782
rect 35808 5296 35860 5302
rect 35912 5284 35940 6326
rect 36636 6248 36688 6254
rect 36636 6190 36688 6196
rect 35860 5256 35940 5284
rect 35808 5238 35860 5244
rect 33232 5160 33284 5166
rect 35072 5160 35124 5166
rect 33232 5102 33284 5108
rect 34900 5108 35072 5114
rect 34900 5102 35124 5108
rect 34900 5086 35112 5102
rect 35256 5092 35308 5098
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 33152 4690 33180 4762
rect 33140 4684 33192 4690
rect 33140 4626 33192 4632
rect 34428 4276 34480 4282
rect 34428 4218 34480 4224
rect 34440 4026 34468 4218
rect 34900 4078 34928 5086
rect 35256 5034 35308 5040
rect 35268 4554 35296 5034
rect 36648 5030 36676 6190
rect 36740 5710 36768 6394
rect 37740 6112 37792 6118
rect 37740 6054 37792 6060
rect 37070 6012 37378 6021
rect 37070 6010 37076 6012
rect 37132 6010 37156 6012
rect 37212 6010 37236 6012
rect 37292 6010 37316 6012
rect 37372 6010 37378 6012
rect 37132 5958 37134 6010
rect 37314 5958 37316 6010
rect 37070 5956 37076 5958
rect 37132 5956 37156 5958
rect 37212 5956 37236 5958
rect 37292 5956 37316 5958
rect 37372 5956 37378 5958
rect 37070 5947 37378 5956
rect 36728 5704 36780 5710
rect 36728 5646 36780 5652
rect 37556 5636 37608 5642
rect 37556 5578 37608 5584
rect 37568 5370 37596 5578
rect 37556 5364 37608 5370
rect 37556 5306 37608 5312
rect 37648 5228 37700 5234
rect 37648 5170 37700 5176
rect 36636 5024 36688 5030
rect 36636 4966 36688 4972
rect 37556 5024 37608 5030
rect 37556 4966 37608 4972
rect 35256 4548 35308 4554
rect 35256 4490 35308 4496
rect 35268 4282 35296 4490
rect 35256 4276 35308 4282
rect 35256 4218 35308 4224
rect 34888 4072 34940 4078
rect 34440 4010 34560 4026
rect 34888 4014 34940 4020
rect 34440 4004 34572 4010
rect 34440 3998 34520 4004
rect 34520 3946 34572 3952
rect 34428 3936 34480 3942
rect 34428 3878 34480 3884
rect 34440 3738 34468 3878
rect 34428 3732 34480 3738
rect 34428 3674 34480 3680
rect 34900 3652 34928 4014
rect 35072 3664 35124 3670
rect 34900 3624 35072 3652
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 34900 3058 34928 3624
rect 35268 3652 35296 4218
rect 36648 4078 36676 4966
rect 37070 4924 37378 4933
rect 37070 4922 37076 4924
rect 37132 4922 37156 4924
rect 37212 4922 37236 4924
rect 37292 4922 37316 4924
rect 37372 4922 37378 4924
rect 37132 4870 37134 4922
rect 37314 4870 37316 4922
rect 37070 4868 37076 4870
rect 37132 4868 37156 4870
rect 37212 4868 37236 4870
rect 37292 4868 37316 4870
rect 37372 4868 37378 4870
rect 37070 4859 37378 4868
rect 37568 4078 37596 4966
rect 37660 4826 37688 5170
rect 37752 5166 37780 6054
rect 37740 5160 37792 5166
rect 37740 5102 37792 5108
rect 37648 4820 37700 4826
rect 37648 4762 37700 4768
rect 37740 4548 37792 4554
rect 37740 4490 37792 4496
rect 37752 4146 37780 4490
rect 37740 4140 37792 4146
rect 37740 4082 37792 4088
rect 36636 4072 36688 4078
rect 36636 4014 36688 4020
rect 37556 4072 37608 4078
rect 37556 4014 37608 4020
rect 37070 3836 37378 3845
rect 37070 3834 37076 3836
rect 37132 3834 37156 3836
rect 37212 3834 37236 3836
rect 37292 3834 37316 3836
rect 37372 3834 37378 3836
rect 37132 3782 37134 3834
rect 37314 3782 37316 3834
rect 37070 3780 37076 3782
rect 37132 3780 37156 3782
rect 37212 3780 37236 3782
rect 37292 3780 37316 3782
rect 37372 3780 37378 3782
rect 37070 3771 37378 3780
rect 35072 3606 35124 3612
rect 35176 3624 35296 3652
rect 35176 3466 35204 3624
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 29184 2984 29236 2990
rect 29184 2926 29236 2932
rect 29552 2916 29604 2922
rect 29552 2858 29604 2864
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19720 2446 19748 2790
rect 22622 2748 22930 2757
rect 22622 2746 22628 2748
rect 22684 2746 22708 2748
rect 22764 2746 22788 2748
rect 22844 2746 22868 2748
rect 22924 2746 22930 2748
rect 22684 2694 22686 2746
rect 22866 2694 22868 2746
rect 22622 2692 22628 2694
rect 22684 2692 22708 2694
rect 22764 2692 22788 2694
rect 22844 2692 22868 2694
rect 22924 2692 22930 2694
rect 22622 2683 22930 2692
rect 29564 2446 29592 2858
rect 33784 2848 33836 2854
rect 33784 2790 33836 2796
rect 33796 2446 33824 2790
rect 37070 2748 37378 2757
rect 37070 2746 37076 2748
rect 37132 2746 37156 2748
rect 37212 2746 37236 2748
rect 37292 2746 37316 2748
rect 37372 2746 37378 2748
rect 37132 2694 37134 2746
rect 37314 2694 37316 2746
rect 37070 2692 37076 2694
rect 37132 2692 37156 2694
rect 37212 2692 37236 2694
rect 37292 2692 37316 2694
rect 37372 2692 37378 2694
rect 37070 2683 37378 2692
rect 37844 2650 37872 11308
rect 37936 11014 37964 11784
rect 38212 11558 38240 13126
rect 38292 12096 38344 12102
rect 38292 12038 38344 12044
rect 38304 11558 38332 12038
rect 38200 11552 38252 11558
rect 38200 11494 38252 11500
rect 38292 11552 38344 11558
rect 38292 11494 38344 11500
rect 38108 11144 38160 11150
rect 38106 11112 38108 11121
rect 38160 11112 38162 11121
rect 38212 11082 38240 11494
rect 38106 11047 38162 11056
rect 38200 11076 38252 11082
rect 37924 11008 37976 11014
rect 37924 10950 37976 10956
rect 37936 10674 37964 10950
rect 37924 10668 37976 10674
rect 37924 10610 37976 10616
rect 38120 9926 38148 11047
rect 38200 11018 38252 11024
rect 38212 9994 38240 11018
rect 38200 9988 38252 9994
rect 38200 9930 38252 9936
rect 38108 9920 38160 9926
rect 38108 9862 38160 9868
rect 38212 9042 38240 9930
rect 38396 9654 38424 15370
rect 38672 14482 38700 15506
rect 38948 15502 38976 17682
rect 39120 17604 39172 17610
rect 39120 17546 39172 17552
rect 39028 16992 39080 16998
rect 39028 16934 39080 16940
rect 39040 16114 39068 16934
rect 39028 16108 39080 16114
rect 39028 16050 39080 16056
rect 39028 15972 39080 15978
rect 39028 15914 39080 15920
rect 38936 15496 38988 15502
rect 38936 15438 38988 15444
rect 38752 15360 38804 15366
rect 38752 15302 38804 15308
rect 38764 15094 38792 15302
rect 38752 15088 38804 15094
rect 38752 15030 38804 15036
rect 39040 15026 39068 15914
rect 39132 15745 39160 17546
rect 39408 16250 39436 19722
rect 40144 18834 40172 20198
rect 40328 19514 40356 20402
rect 40316 19508 40368 19514
rect 40316 19450 40368 19456
rect 40132 18828 40184 18834
rect 40132 18770 40184 18776
rect 39488 18760 39540 18766
rect 39488 18702 39540 18708
rect 39500 18086 39528 18702
rect 39488 18080 39540 18086
rect 39488 18022 39540 18028
rect 39500 17202 39528 18022
rect 40328 17678 40356 19450
rect 40316 17672 40368 17678
rect 40316 17614 40368 17620
rect 39488 17196 39540 17202
rect 39488 17138 39540 17144
rect 39764 17128 39816 17134
rect 39764 17070 39816 17076
rect 39776 16794 39804 17070
rect 39764 16788 39816 16794
rect 39764 16730 39816 16736
rect 39396 16244 39448 16250
rect 39396 16186 39448 16192
rect 39672 16108 39724 16114
rect 39672 16050 39724 16056
rect 39118 15736 39174 15745
rect 39118 15671 39174 15680
rect 39684 15638 39712 16050
rect 39672 15632 39724 15638
rect 39672 15574 39724 15580
rect 39948 15564 40000 15570
rect 39948 15506 40000 15512
rect 39960 15162 39988 15506
rect 39948 15156 40000 15162
rect 39948 15098 40000 15104
rect 39028 15020 39080 15026
rect 39028 14962 39080 14968
rect 38660 14476 38712 14482
rect 38660 14418 38712 14424
rect 39304 14340 39356 14346
rect 39304 14282 39356 14288
rect 39316 13870 39344 14282
rect 39304 13864 39356 13870
rect 39304 13806 39356 13812
rect 39396 13864 39448 13870
rect 39396 13806 39448 13812
rect 39408 12986 39436 13806
rect 39960 13530 39988 15098
rect 40132 15020 40184 15026
rect 40132 14962 40184 14968
rect 40144 14278 40172 14962
rect 40500 14952 40552 14958
rect 40500 14894 40552 14900
rect 40132 14272 40184 14278
rect 40132 14214 40184 14220
rect 40040 13932 40092 13938
rect 40040 13874 40092 13880
rect 40052 13530 40080 13874
rect 39948 13524 40000 13530
rect 39948 13466 40000 13472
rect 40040 13524 40092 13530
rect 40040 13466 40092 13472
rect 39396 12980 39448 12986
rect 39396 12922 39448 12928
rect 39408 12850 39436 12922
rect 39396 12844 39448 12850
rect 39396 12786 39448 12792
rect 40144 12782 40172 14214
rect 40512 13326 40540 14894
rect 40604 14414 40632 20402
rect 41236 20256 41288 20262
rect 41236 20198 41288 20204
rect 40684 20052 40736 20058
rect 40684 19994 40736 20000
rect 40696 16658 40724 19994
rect 40868 19916 40920 19922
rect 40868 19858 40920 19864
rect 40880 18290 40908 19858
rect 41052 19440 41104 19446
rect 41052 19382 41104 19388
rect 41064 18426 41092 19382
rect 41248 18766 41276 20198
rect 41340 19922 41368 20742
rect 41788 20256 41840 20262
rect 41788 20198 41840 20204
rect 41696 19984 41748 19990
rect 41800 19961 41828 20198
rect 41696 19926 41748 19932
rect 41786 19952 41842 19961
rect 41328 19916 41380 19922
rect 41328 19858 41380 19864
rect 41604 19372 41656 19378
rect 41604 19314 41656 19320
rect 41236 18760 41288 18766
rect 41236 18702 41288 18708
rect 41616 18630 41644 19314
rect 41420 18624 41472 18630
rect 41604 18624 41656 18630
rect 41472 18584 41552 18612
rect 41420 18566 41472 18572
rect 41052 18420 41104 18426
rect 41052 18362 41104 18368
rect 40868 18284 40920 18290
rect 40868 18226 40920 18232
rect 40776 17264 40828 17270
rect 40776 17206 40828 17212
rect 40788 16794 40816 17206
rect 40776 16788 40828 16794
rect 40776 16730 40828 16736
rect 40684 16652 40736 16658
rect 40684 16594 40736 16600
rect 40696 15162 40724 16594
rect 40880 15502 40908 18226
rect 41420 18216 41472 18222
rect 41420 18158 41472 18164
rect 41432 18086 41460 18158
rect 41420 18080 41472 18086
rect 41420 18022 41472 18028
rect 41420 17876 41472 17882
rect 41420 17818 41472 17824
rect 41236 17672 41288 17678
rect 41236 17614 41288 17620
rect 40960 17536 41012 17542
rect 41248 17524 41276 17614
rect 41012 17496 41276 17524
rect 40960 17478 41012 17484
rect 41236 16992 41288 16998
rect 41236 16934 41288 16940
rect 41052 16448 41104 16454
rect 41052 16390 41104 16396
rect 41064 16114 41092 16390
rect 41052 16108 41104 16114
rect 41052 16050 41104 16056
rect 41248 16046 41276 16934
rect 41328 16448 41380 16454
rect 41328 16390 41380 16396
rect 41236 16040 41288 16046
rect 41236 15982 41288 15988
rect 40868 15496 40920 15502
rect 40868 15438 40920 15444
rect 40684 15156 40736 15162
rect 40684 15098 40736 15104
rect 41144 15020 41196 15026
rect 41144 14962 41196 14968
rect 41156 14414 41184 14962
rect 40592 14408 40644 14414
rect 40592 14350 40644 14356
rect 40684 14408 40736 14414
rect 40684 14350 40736 14356
rect 41144 14408 41196 14414
rect 41144 14350 41196 14356
rect 40696 14006 40724 14350
rect 40684 14000 40736 14006
rect 40684 13942 40736 13948
rect 40696 13870 40724 13942
rect 40960 13932 41012 13938
rect 41156 13920 41184 14350
rect 41012 13892 41184 13920
rect 40960 13874 41012 13880
rect 40684 13864 40736 13870
rect 40684 13806 40736 13812
rect 40592 13524 40644 13530
rect 40592 13466 40644 13472
rect 40500 13320 40552 13326
rect 40500 13262 40552 13268
rect 40132 12776 40184 12782
rect 40132 12718 40184 12724
rect 38476 12640 38528 12646
rect 38476 12582 38528 12588
rect 40132 12640 40184 12646
rect 40132 12582 40184 12588
rect 38488 12238 38516 12582
rect 38752 12436 38804 12442
rect 38752 12378 38804 12384
rect 38764 12238 38792 12378
rect 39856 12368 39908 12374
rect 39856 12310 39908 12316
rect 39764 12300 39816 12306
rect 39764 12242 39816 12248
rect 38476 12232 38528 12238
rect 38476 12174 38528 12180
rect 38752 12232 38804 12238
rect 38752 12174 38804 12180
rect 39776 12170 39804 12242
rect 39868 12238 39896 12310
rect 40144 12238 40172 12582
rect 40512 12306 40540 13262
rect 40604 12850 40632 13466
rect 40696 13394 40724 13806
rect 40684 13388 40736 13394
rect 40684 13330 40736 13336
rect 40972 13308 41000 13874
rect 41144 13320 41196 13326
rect 40972 13280 41144 13308
rect 40972 12986 41000 13280
rect 41144 13262 41196 13268
rect 40960 12980 41012 12986
rect 40960 12922 41012 12928
rect 40972 12850 41000 12922
rect 40592 12844 40644 12850
rect 40592 12786 40644 12792
rect 40960 12844 41012 12850
rect 40960 12786 41012 12792
rect 40500 12300 40552 12306
rect 40500 12242 40552 12248
rect 41156 12238 41184 13262
rect 41340 13258 41368 16390
rect 41432 15094 41460 17818
rect 41524 16522 41552 18584
rect 41604 18566 41656 18572
rect 41616 17746 41644 18566
rect 41708 18290 41736 19926
rect 41786 19887 41788 19896
rect 41840 19887 41842 19896
rect 41788 19858 41840 19864
rect 41800 19827 41828 19858
rect 41696 18284 41748 18290
rect 41696 18226 41748 18232
rect 41604 17740 41656 17746
rect 41604 17682 41656 17688
rect 41512 16516 41564 16522
rect 41512 16458 41564 16464
rect 41708 16250 41736 18226
rect 41892 17882 41920 22510
rect 42536 22438 42564 22578
rect 42524 22432 42576 22438
rect 42524 22374 42576 22380
rect 42536 22094 42564 22374
rect 42536 22066 42656 22094
rect 42628 21486 42656 22066
rect 43444 22024 43496 22030
rect 43444 21966 43496 21972
rect 42616 21480 42668 21486
rect 42616 21422 42668 21428
rect 42708 21480 42760 21486
rect 42708 21422 42760 21428
rect 42628 21078 42656 21422
rect 42616 21072 42668 21078
rect 42616 21014 42668 21020
rect 42720 21010 42748 21422
rect 43456 21350 43484 21966
rect 43628 21412 43680 21418
rect 43628 21354 43680 21360
rect 43444 21344 43496 21350
rect 43444 21286 43496 21292
rect 42984 21140 43036 21146
rect 42984 21082 43036 21088
rect 42708 21004 42760 21010
rect 42708 20946 42760 20952
rect 42432 20868 42484 20874
rect 42432 20810 42484 20816
rect 42444 20262 42472 20810
rect 42996 20466 43024 21082
rect 43352 20528 43404 20534
rect 43352 20470 43404 20476
rect 42984 20460 43036 20466
rect 42984 20402 43036 20408
rect 42432 20256 42484 20262
rect 42432 20198 42484 20204
rect 42064 19848 42116 19854
rect 42064 19790 42116 19796
rect 42076 18358 42104 19790
rect 42156 19712 42208 19718
rect 42156 19654 42208 19660
rect 42168 19514 42196 19654
rect 42156 19508 42208 19514
rect 42156 19450 42208 19456
rect 42444 18766 42472 20198
rect 42616 20052 42668 20058
rect 42616 19994 42668 20000
rect 42628 19378 42656 19994
rect 42616 19372 42668 19378
rect 42616 19314 42668 19320
rect 42432 18760 42484 18766
rect 42432 18702 42484 18708
rect 42800 18624 42852 18630
rect 42800 18566 42852 18572
rect 42352 18414 42656 18442
rect 42064 18352 42116 18358
rect 42064 18294 42116 18300
rect 41880 17876 41932 17882
rect 41880 17818 41932 17824
rect 42076 17678 42104 18294
rect 42352 18222 42380 18414
rect 42524 18352 42576 18358
rect 42524 18294 42576 18300
rect 42340 18216 42392 18222
rect 42536 18170 42564 18294
rect 42628 18290 42656 18414
rect 42616 18284 42668 18290
rect 42616 18226 42668 18232
rect 42340 18158 42392 18164
rect 42444 18154 42564 18170
rect 42432 18148 42564 18154
rect 42484 18142 42564 18148
rect 42432 18090 42484 18096
rect 42536 17882 42564 18142
rect 42524 17876 42576 17882
rect 42524 17818 42576 17824
rect 42064 17672 42116 17678
rect 42064 17614 42116 17620
rect 41788 17536 41840 17542
rect 41788 17478 41840 17484
rect 41800 17202 41828 17478
rect 41788 17196 41840 17202
rect 41788 17138 41840 17144
rect 41800 16726 41828 17138
rect 41788 16720 41840 16726
rect 41788 16662 41840 16668
rect 42628 16658 42656 18226
rect 42812 17610 42840 18566
rect 42996 18086 43024 20402
rect 43076 20256 43128 20262
rect 43076 20198 43128 20204
rect 43088 19378 43116 20198
rect 43260 19916 43312 19922
rect 43260 19858 43312 19864
rect 43272 19514 43300 19858
rect 43260 19508 43312 19514
rect 43260 19450 43312 19456
rect 43076 19372 43128 19378
rect 43076 19314 43128 19320
rect 43088 18834 43116 19314
rect 43076 18828 43128 18834
rect 43076 18770 43128 18776
rect 43364 18290 43392 20470
rect 43352 18284 43404 18290
rect 43352 18226 43404 18232
rect 43364 18193 43392 18226
rect 43350 18184 43406 18193
rect 43350 18119 43406 18128
rect 42984 18080 43036 18086
rect 42984 18022 43036 18028
rect 42892 17808 42944 17814
rect 42892 17750 42944 17756
rect 42800 17604 42852 17610
rect 42800 17546 42852 17552
rect 42812 16794 42840 17546
rect 42904 17134 42932 17750
rect 42892 17128 42944 17134
rect 42892 17070 42944 17076
rect 42800 16788 42852 16794
rect 42800 16730 42852 16736
rect 43168 16720 43220 16726
rect 43456 16674 43484 21286
rect 43640 21010 43668 21354
rect 43628 21004 43680 21010
rect 43628 20946 43680 20952
rect 43628 20392 43680 20398
rect 43628 20334 43680 20340
rect 43640 20058 43668 20334
rect 43628 20052 43680 20058
rect 43628 19994 43680 20000
rect 43536 19848 43588 19854
rect 43536 19790 43588 19796
rect 43548 18766 43576 19790
rect 43536 18760 43588 18766
rect 43536 18702 43588 18708
rect 43548 17066 43576 18702
rect 43812 18148 43864 18154
rect 43812 18090 43864 18096
rect 43824 17746 43852 18090
rect 43812 17740 43864 17746
rect 43812 17682 43864 17688
rect 43536 17060 43588 17066
rect 43536 17002 43588 17008
rect 43220 16668 43668 16674
rect 43168 16662 43668 16668
rect 42616 16652 42668 16658
rect 43180 16646 43668 16662
rect 42616 16594 42668 16600
rect 41696 16244 41748 16250
rect 41696 16186 41748 16192
rect 42064 16176 42116 16182
rect 42064 16118 42116 16124
rect 41880 16040 41932 16046
rect 41880 15982 41932 15988
rect 41602 15736 41658 15745
rect 41892 15706 41920 15982
rect 41602 15671 41658 15680
rect 41880 15700 41932 15706
rect 41420 15088 41472 15094
rect 41420 15030 41472 15036
rect 41420 14952 41472 14958
rect 41420 14894 41472 14900
rect 41432 14414 41460 14894
rect 41420 14408 41472 14414
rect 41420 14350 41472 14356
rect 41328 13252 41380 13258
rect 41328 13194 41380 13200
rect 41340 12434 41368 13194
rect 41512 12708 41564 12714
rect 41512 12650 41564 12656
rect 41524 12442 41552 12650
rect 41248 12406 41368 12434
rect 41512 12436 41564 12442
rect 39856 12232 39908 12238
rect 39856 12174 39908 12180
rect 40132 12232 40184 12238
rect 40132 12174 40184 12180
rect 41144 12232 41196 12238
rect 41144 12174 41196 12180
rect 39580 12164 39632 12170
rect 39580 12106 39632 12112
rect 39764 12164 39816 12170
rect 39764 12106 39816 12112
rect 38568 11824 38620 11830
rect 38488 11784 38568 11812
rect 38488 11694 38516 11784
rect 38568 11766 38620 11772
rect 39592 11694 39620 12106
rect 40040 12096 40092 12102
rect 39960 12056 40040 12084
rect 38476 11688 38528 11694
rect 38476 11630 38528 11636
rect 38844 11688 38896 11694
rect 38844 11630 38896 11636
rect 39580 11688 39632 11694
rect 39580 11630 39632 11636
rect 38488 11150 38516 11630
rect 38856 11354 38884 11630
rect 38844 11348 38896 11354
rect 38844 11290 38896 11296
rect 39960 11218 39988 12056
rect 40040 12038 40092 12044
rect 40144 11286 40172 12174
rect 40684 11824 40736 11830
rect 40684 11766 40736 11772
rect 40592 11756 40644 11762
rect 40592 11698 40644 11704
rect 40224 11620 40276 11626
rect 40224 11562 40276 11568
rect 40132 11280 40184 11286
rect 40132 11222 40184 11228
rect 39948 11212 40000 11218
rect 39948 11154 40000 11160
rect 38476 11144 38528 11150
rect 38476 11086 38528 11092
rect 40040 11144 40092 11150
rect 40040 11086 40092 11092
rect 38476 10804 38528 10810
rect 38476 10746 38528 10752
rect 38488 10713 38516 10746
rect 38936 10736 38988 10742
rect 38474 10704 38530 10713
rect 38936 10678 38988 10684
rect 39212 10736 39264 10742
rect 39212 10678 39264 10684
rect 38474 10639 38530 10648
rect 38660 10124 38712 10130
rect 38660 10066 38712 10072
rect 38672 10033 38700 10066
rect 38658 10024 38714 10033
rect 38476 9988 38528 9994
rect 38658 9959 38714 9968
rect 38476 9930 38528 9936
rect 38384 9648 38436 9654
rect 38384 9590 38436 9596
rect 38200 9036 38252 9042
rect 38200 8978 38252 8984
rect 38016 8968 38068 8974
rect 38016 8910 38068 8916
rect 38292 8968 38344 8974
rect 38292 8910 38344 8916
rect 38028 7818 38056 8910
rect 38016 7812 38068 7818
rect 38016 7754 38068 7760
rect 38304 6905 38332 8910
rect 38488 8634 38516 9930
rect 38844 9512 38896 9518
rect 38844 9454 38896 9460
rect 38568 9172 38620 9178
rect 38568 9114 38620 9120
rect 38476 8628 38528 8634
rect 38476 8570 38528 8576
rect 38580 8498 38608 9114
rect 38660 9104 38712 9110
rect 38752 9104 38804 9110
rect 38712 9064 38752 9092
rect 38660 9046 38712 9052
rect 38752 9046 38804 9052
rect 38856 8974 38884 9454
rect 38948 9382 38976 10678
rect 39120 10056 39172 10062
rect 39120 9998 39172 10004
rect 38936 9376 38988 9382
rect 38936 9318 38988 9324
rect 38660 8968 38712 8974
rect 38660 8910 38712 8916
rect 38844 8968 38896 8974
rect 38844 8910 38896 8916
rect 38672 8673 38700 8910
rect 38658 8664 38714 8673
rect 38658 8599 38714 8608
rect 38568 8492 38620 8498
rect 38568 8434 38620 8440
rect 38384 8424 38436 8430
rect 38384 8366 38436 8372
rect 38396 7546 38424 8366
rect 38476 8356 38528 8362
rect 38476 8298 38528 8304
rect 38488 7954 38516 8298
rect 38476 7948 38528 7954
rect 38476 7890 38528 7896
rect 38476 7812 38528 7818
rect 38476 7754 38528 7760
rect 38488 7546 38516 7754
rect 38384 7540 38436 7546
rect 38384 7482 38436 7488
rect 38476 7540 38528 7546
rect 38476 7482 38528 7488
rect 38290 6896 38346 6905
rect 38290 6831 38346 6840
rect 38016 6724 38068 6730
rect 38016 6666 38068 6672
rect 37924 6316 37976 6322
rect 37924 6258 37976 6264
rect 37936 5914 37964 6258
rect 37924 5908 37976 5914
rect 37924 5850 37976 5856
rect 38028 5642 38056 6666
rect 38200 6384 38252 6390
rect 38200 6326 38252 6332
rect 38016 5636 38068 5642
rect 38016 5578 38068 5584
rect 38028 3126 38056 5578
rect 38108 5228 38160 5234
rect 38108 5170 38160 5176
rect 38120 4622 38148 5170
rect 38212 4690 38240 6326
rect 38304 5166 38332 6831
rect 38488 6798 38516 7482
rect 38580 7342 38608 8434
rect 38568 7336 38620 7342
rect 38568 7278 38620 7284
rect 38856 6798 38884 8910
rect 38476 6792 38528 6798
rect 38476 6734 38528 6740
rect 38844 6792 38896 6798
rect 38844 6734 38896 6740
rect 38752 6316 38804 6322
rect 38752 6258 38804 6264
rect 38292 5160 38344 5166
rect 38292 5102 38344 5108
rect 38200 4684 38252 4690
rect 38200 4626 38252 4632
rect 38764 4622 38792 6258
rect 38948 5574 38976 9318
rect 39132 9042 39160 9998
rect 39120 9036 39172 9042
rect 39120 8978 39172 8984
rect 39028 8968 39080 8974
rect 39028 8910 39080 8916
rect 39040 7993 39068 8910
rect 39120 8832 39172 8838
rect 39120 8774 39172 8780
rect 39132 8566 39160 8774
rect 39120 8560 39172 8566
rect 39120 8502 39172 8508
rect 39026 7984 39082 7993
rect 39026 7919 39082 7928
rect 39040 6866 39068 7919
rect 39028 6860 39080 6866
rect 39028 6802 39080 6808
rect 39132 6798 39160 8502
rect 39224 7342 39252 10678
rect 40052 10538 40080 11086
rect 40040 10532 40092 10538
rect 40040 10474 40092 10480
rect 39948 10464 40000 10470
rect 39948 10406 40000 10412
rect 39304 10056 39356 10062
rect 39304 9998 39356 10004
rect 39316 9450 39344 9998
rect 39304 9444 39356 9450
rect 39304 9386 39356 9392
rect 39316 8906 39344 9386
rect 39764 9376 39816 9382
rect 39764 9318 39816 9324
rect 39304 8900 39356 8906
rect 39304 8842 39356 8848
rect 39316 8566 39344 8842
rect 39304 8560 39356 8566
rect 39776 8537 39804 9318
rect 39960 8634 39988 10406
rect 40052 10130 40080 10474
rect 40236 10470 40264 11562
rect 40316 10668 40368 10674
rect 40316 10610 40368 10616
rect 40224 10464 40276 10470
rect 40224 10406 40276 10412
rect 40236 10130 40264 10406
rect 40040 10124 40092 10130
rect 40040 10066 40092 10072
rect 40224 10124 40276 10130
rect 40224 10066 40276 10072
rect 40052 9654 40080 10066
rect 40132 9920 40184 9926
rect 40132 9862 40184 9868
rect 40144 9722 40172 9862
rect 40132 9716 40184 9722
rect 40132 9658 40184 9664
rect 40040 9648 40092 9654
rect 40040 9590 40092 9596
rect 40052 8974 40080 9590
rect 40040 8968 40092 8974
rect 40040 8910 40092 8916
rect 39948 8628 40000 8634
rect 39948 8570 40000 8576
rect 39304 8502 39356 8508
rect 39762 8528 39818 8537
rect 39762 8463 39818 8472
rect 39856 8492 39908 8498
rect 39856 8434 39908 8440
rect 39672 8424 39724 8430
rect 39868 8401 39896 8434
rect 39948 8424 40000 8430
rect 39672 8366 39724 8372
rect 39854 8392 39910 8401
rect 39684 8265 39712 8366
rect 39764 8356 39816 8362
rect 39948 8366 40000 8372
rect 39854 8327 39910 8336
rect 39764 8298 39816 8304
rect 39670 8256 39726 8265
rect 39670 8191 39726 8200
rect 39776 7478 39804 8298
rect 39868 8022 39896 8327
rect 39960 8294 39988 8366
rect 39948 8288 40000 8294
rect 39948 8230 40000 8236
rect 40236 8090 40264 10066
rect 40328 8974 40356 10610
rect 40604 10266 40632 11698
rect 40592 10260 40644 10266
rect 40592 10202 40644 10208
rect 40316 8968 40368 8974
rect 40368 8928 40540 8956
rect 40316 8910 40368 8916
rect 40512 8294 40540 8928
rect 40408 8288 40460 8294
rect 40408 8230 40460 8236
rect 40500 8288 40552 8294
rect 40500 8230 40552 8236
rect 40224 8084 40276 8090
rect 40224 8026 40276 8032
rect 39856 8016 39908 8022
rect 39856 7958 39908 7964
rect 39764 7472 39816 7478
rect 39764 7414 39816 7420
rect 39212 7336 39264 7342
rect 39212 7278 39264 7284
rect 39868 6866 39896 7958
rect 40040 7948 40092 7954
rect 40040 7890 40092 7896
rect 40052 7410 40080 7890
rect 40420 7818 40448 8230
rect 40408 7812 40460 7818
rect 40408 7754 40460 7760
rect 40408 7472 40460 7478
rect 40408 7414 40460 7420
rect 40040 7404 40092 7410
rect 40040 7346 40092 7352
rect 39856 6860 39908 6866
rect 39856 6802 39908 6808
rect 39120 6792 39172 6798
rect 39120 6734 39172 6740
rect 39868 6322 39896 6802
rect 39856 6316 39908 6322
rect 39856 6258 39908 6264
rect 39028 6112 39080 6118
rect 39028 6054 39080 6060
rect 39040 5846 39068 6054
rect 39028 5840 39080 5846
rect 39028 5782 39080 5788
rect 38936 5568 38988 5574
rect 38936 5510 38988 5516
rect 38948 5302 38976 5510
rect 38936 5296 38988 5302
rect 38936 5238 38988 5244
rect 39040 4690 39068 5782
rect 39948 5568 40000 5574
rect 39948 5510 40000 5516
rect 39856 5092 39908 5098
rect 39856 5034 39908 5040
rect 39028 4684 39080 4690
rect 39028 4626 39080 4632
rect 39868 4622 39896 5034
rect 39960 5030 39988 5510
rect 40052 5370 40080 7346
rect 40420 6798 40448 7414
rect 40408 6792 40460 6798
rect 40408 6734 40460 6740
rect 40696 6730 40724 11766
rect 40960 11756 41012 11762
rect 40960 11698 41012 11704
rect 40972 11286 41000 11698
rect 40776 11280 40828 11286
rect 40776 11222 40828 11228
rect 40960 11280 41012 11286
rect 40960 11222 41012 11228
rect 40788 10266 40816 11222
rect 40972 10810 41000 11222
rect 41248 11218 41276 12406
rect 41512 12378 41564 12384
rect 41236 11212 41288 11218
rect 41236 11154 41288 11160
rect 40960 10804 41012 10810
rect 40960 10746 41012 10752
rect 40776 10260 40828 10266
rect 40776 10202 40828 10208
rect 40972 9602 41000 10746
rect 41144 10532 41196 10538
rect 41144 10474 41196 10480
rect 41156 9926 41184 10474
rect 41248 10130 41276 11154
rect 41420 10192 41472 10198
rect 41420 10134 41472 10140
rect 41236 10124 41288 10130
rect 41236 10066 41288 10072
rect 41144 9920 41196 9926
rect 41144 9862 41196 9868
rect 41236 9920 41288 9926
rect 41236 9862 41288 9868
rect 40880 9574 41000 9602
rect 40880 9382 40908 9574
rect 40960 9512 41012 9518
rect 40960 9454 41012 9460
rect 40868 9376 40920 9382
rect 40868 9318 40920 9324
rect 40880 9178 40908 9318
rect 40868 9172 40920 9178
rect 40868 9114 40920 9120
rect 40866 8664 40922 8673
rect 40972 8634 41000 9454
rect 41052 9376 41104 9382
rect 41052 9318 41104 9324
rect 40866 8599 40922 8608
rect 40960 8628 41012 8634
rect 40880 8412 40908 8599
rect 40960 8570 41012 8576
rect 40960 8424 41012 8430
rect 40880 8384 40960 8412
rect 41064 8412 41092 9318
rect 41012 8384 41092 8412
rect 40960 8366 41012 8372
rect 41156 7546 41184 9862
rect 41248 9654 41276 9862
rect 41236 9648 41288 9654
rect 41236 9590 41288 9596
rect 41328 9580 41380 9586
rect 41328 9522 41380 9528
rect 41340 9178 41368 9522
rect 41328 9172 41380 9178
rect 41328 9114 41380 9120
rect 41432 8514 41460 10134
rect 41432 8486 41552 8514
rect 41616 8498 41644 15671
rect 41880 15642 41932 15648
rect 41880 15428 41932 15434
rect 41880 15370 41932 15376
rect 41892 15094 41920 15370
rect 41880 15088 41932 15094
rect 41880 15030 41932 15036
rect 41788 15020 41840 15026
rect 41788 14962 41840 14968
rect 41696 14408 41748 14414
rect 41696 14350 41748 14356
rect 41708 14074 41736 14350
rect 41800 14346 41828 14962
rect 41788 14340 41840 14346
rect 41788 14282 41840 14288
rect 41696 14068 41748 14074
rect 41696 14010 41748 14016
rect 41708 13938 41736 14010
rect 41696 13932 41748 13938
rect 41696 13874 41748 13880
rect 41708 13326 41736 13874
rect 41696 13320 41748 13326
rect 41696 13262 41748 13268
rect 41708 12986 41736 13262
rect 41696 12980 41748 12986
rect 41696 12922 41748 12928
rect 41800 12434 41828 14282
rect 42076 14278 42104 16118
rect 42628 14958 42656 16594
rect 42616 14952 42668 14958
rect 42616 14894 42668 14900
rect 42892 14952 42944 14958
rect 42892 14894 42944 14900
rect 42524 14544 42576 14550
rect 42576 14504 42656 14532
rect 42524 14486 42576 14492
rect 42524 14340 42576 14346
rect 42524 14282 42576 14288
rect 42064 14272 42116 14278
rect 42064 14214 42116 14220
rect 42536 14006 42564 14282
rect 42524 14000 42576 14006
rect 42524 13942 42576 13948
rect 42156 13728 42208 13734
rect 42156 13670 42208 13676
rect 42168 13258 42196 13670
rect 42628 13530 42656 14504
rect 42904 14414 42932 14894
rect 42984 14816 43036 14822
rect 42984 14758 43036 14764
rect 42892 14408 42944 14414
rect 42720 14368 42892 14396
rect 42720 13938 42748 14368
rect 42892 14350 42944 14356
rect 42996 14278 43024 14758
rect 43536 14408 43588 14414
rect 43536 14350 43588 14356
rect 42984 14272 43036 14278
rect 42984 14214 43036 14220
rect 43444 14000 43496 14006
rect 43444 13942 43496 13948
rect 42708 13932 42760 13938
rect 42760 13892 42840 13920
rect 42708 13874 42760 13880
rect 42616 13524 42668 13530
rect 42616 13466 42668 13472
rect 42628 13394 42656 13466
rect 42616 13388 42668 13394
rect 42616 13330 42668 13336
rect 42812 13326 42840 13892
rect 42800 13320 42852 13326
rect 42800 13262 42852 13268
rect 42156 13252 42208 13258
rect 42156 13194 42208 13200
rect 42168 12782 42196 13194
rect 42156 12776 42208 12782
rect 42156 12718 42208 12724
rect 42168 12442 42196 12718
rect 42156 12436 42208 12442
rect 41800 12406 42012 12434
rect 41984 12238 42012 12406
rect 42076 12406 42156 12434
rect 41972 12232 42024 12238
rect 41972 12174 42024 12180
rect 41984 11898 42012 12174
rect 41972 11892 42024 11898
rect 41972 11834 42024 11840
rect 41420 8356 41472 8362
rect 41420 8298 41472 8304
rect 41328 8288 41380 8294
rect 41328 8230 41380 8236
rect 41144 7540 41196 7546
rect 41144 7482 41196 7488
rect 41340 7410 41368 8230
rect 41328 7404 41380 7410
rect 41328 7346 41380 7352
rect 40684 6724 40736 6730
rect 40684 6666 40736 6672
rect 40408 6656 40460 6662
rect 40408 6598 40460 6604
rect 40132 6112 40184 6118
rect 40132 6054 40184 6060
rect 40040 5364 40092 5370
rect 40040 5306 40092 5312
rect 39948 5024 40000 5030
rect 39948 4966 40000 4972
rect 39960 4826 39988 4966
rect 39948 4820 40000 4826
rect 39948 4762 40000 4768
rect 38108 4616 38160 4622
rect 38108 4558 38160 4564
rect 38752 4616 38804 4622
rect 38752 4558 38804 4564
rect 39856 4616 39908 4622
rect 39856 4558 39908 4564
rect 40144 3466 40172 6054
rect 40224 5704 40276 5710
rect 40224 5646 40276 5652
rect 40236 5234 40264 5646
rect 40316 5364 40368 5370
rect 40316 5306 40368 5312
rect 40224 5228 40276 5234
rect 40224 5170 40276 5176
rect 40328 4078 40356 5306
rect 40420 4214 40448 6598
rect 40696 6254 40724 6666
rect 40684 6248 40736 6254
rect 40684 6190 40736 6196
rect 40592 6180 40644 6186
rect 40592 6122 40644 6128
rect 40604 5778 40632 6122
rect 40592 5772 40644 5778
rect 40592 5714 40644 5720
rect 40604 4282 40632 5714
rect 41328 4548 41380 4554
rect 41328 4490 41380 4496
rect 40592 4276 40644 4282
rect 40592 4218 40644 4224
rect 41340 4214 41368 4490
rect 40408 4208 40460 4214
rect 40408 4150 40460 4156
rect 41328 4208 41380 4214
rect 41328 4150 41380 4156
rect 40316 4072 40368 4078
rect 40316 4014 40368 4020
rect 40328 3618 40356 4014
rect 40236 3602 40356 3618
rect 40224 3596 40356 3602
rect 40276 3590 40356 3596
rect 40224 3538 40276 3544
rect 40420 3466 40448 4150
rect 40132 3460 40184 3466
rect 40132 3402 40184 3408
rect 40408 3460 40460 3466
rect 40408 3402 40460 3408
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 41236 3120 41288 3126
rect 41236 3062 41288 3068
rect 41248 2650 41276 3062
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 41236 2644 41288 2650
rect 41236 2586 41288 2592
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 41432 2378 41460 8298
rect 41524 6322 41552 8486
rect 41604 8492 41656 8498
rect 41604 8434 41656 8440
rect 41696 7812 41748 7818
rect 41696 7754 41748 7760
rect 41708 7478 41736 7754
rect 41696 7472 41748 7478
rect 41696 7414 41748 7420
rect 41880 6656 41932 6662
rect 41880 6598 41932 6604
rect 41892 6458 41920 6598
rect 41880 6452 41932 6458
rect 41880 6394 41932 6400
rect 41788 6384 41840 6390
rect 41788 6326 41840 6332
rect 41512 6316 41564 6322
rect 41512 6258 41564 6264
rect 41524 6202 41552 6258
rect 41524 6174 41644 6202
rect 41512 5704 41564 5710
rect 41512 5646 41564 5652
rect 41524 5370 41552 5646
rect 41512 5364 41564 5370
rect 41512 5306 41564 5312
rect 41616 5302 41644 6174
rect 41800 5302 41828 6326
rect 41604 5296 41656 5302
rect 41604 5238 41656 5244
rect 41788 5296 41840 5302
rect 41788 5238 41840 5244
rect 41512 5228 41564 5234
rect 41512 5170 41564 5176
rect 41524 4826 41552 5170
rect 41512 4820 41564 4826
rect 41512 4762 41564 4768
rect 41616 4758 41644 5238
rect 41604 4752 41656 4758
rect 41604 4694 41656 4700
rect 41800 3670 41828 5238
rect 42076 4593 42104 12406
rect 42156 12378 42208 12384
rect 42432 12164 42484 12170
rect 42432 12106 42484 12112
rect 42156 12096 42208 12102
rect 42156 12038 42208 12044
rect 42168 11082 42196 12038
rect 42444 11762 42472 12106
rect 42432 11756 42484 11762
rect 42484 11716 42564 11744
rect 42432 11698 42484 11704
rect 42432 11552 42484 11558
rect 42432 11494 42484 11500
rect 42444 11082 42472 11494
rect 42156 11076 42208 11082
rect 42156 11018 42208 11024
rect 42432 11076 42484 11082
rect 42432 11018 42484 11024
rect 42340 11008 42392 11014
rect 42340 10950 42392 10956
rect 42352 10810 42380 10950
rect 42340 10804 42392 10810
rect 42340 10746 42392 10752
rect 42536 10674 42564 11716
rect 43456 11694 43484 13942
rect 43548 13802 43576 14350
rect 43536 13796 43588 13802
rect 43536 13738 43588 13744
rect 43548 13326 43576 13738
rect 43536 13320 43588 13326
rect 43536 13262 43588 13268
rect 43548 12850 43576 13262
rect 43536 12844 43588 12850
rect 43536 12786 43588 12792
rect 43640 12170 43668 16646
rect 43916 16454 43944 33458
rect 48424 32774 48452 33458
rect 51518 33212 51826 33221
rect 51518 33210 51524 33212
rect 51580 33210 51604 33212
rect 51660 33210 51684 33212
rect 51740 33210 51764 33212
rect 51820 33210 51826 33212
rect 51580 33158 51582 33210
rect 51762 33158 51764 33210
rect 51518 33156 51524 33158
rect 51580 33156 51604 33158
rect 51660 33156 51684 33158
rect 51740 33156 51764 33158
rect 51820 33156 51826 33158
rect 51518 33147 51826 33156
rect 52656 32774 52684 33458
rect 56600 33448 56652 33454
rect 56600 33390 56652 33396
rect 48412 32768 48464 32774
rect 48412 32710 48464 32716
rect 52644 32768 52696 32774
rect 52644 32710 52696 32716
rect 44294 32668 44602 32677
rect 44294 32666 44300 32668
rect 44356 32666 44380 32668
rect 44436 32666 44460 32668
rect 44516 32666 44540 32668
rect 44596 32666 44602 32668
rect 44356 32614 44358 32666
rect 44538 32614 44540 32666
rect 44294 32612 44300 32614
rect 44356 32612 44380 32614
rect 44436 32612 44460 32614
rect 44516 32612 44540 32614
rect 44596 32612 44602 32614
rect 44294 32603 44602 32612
rect 51518 32124 51826 32133
rect 51518 32122 51524 32124
rect 51580 32122 51604 32124
rect 51660 32122 51684 32124
rect 51740 32122 51764 32124
rect 51820 32122 51826 32124
rect 51580 32070 51582 32122
rect 51762 32070 51764 32122
rect 51518 32068 51524 32070
rect 51580 32068 51604 32070
rect 51660 32068 51684 32070
rect 51740 32068 51764 32070
rect 51820 32068 51826 32070
rect 51518 32059 51826 32068
rect 44294 31580 44602 31589
rect 44294 31578 44300 31580
rect 44356 31578 44380 31580
rect 44436 31578 44460 31580
rect 44516 31578 44540 31580
rect 44596 31578 44602 31580
rect 44356 31526 44358 31578
rect 44538 31526 44540 31578
rect 44294 31524 44300 31526
rect 44356 31524 44380 31526
rect 44436 31524 44460 31526
rect 44516 31524 44540 31526
rect 44596 31524 44602 31526
rect 44294 31515 44602 31524
rect 45836 31340 45888 31346
rect 45836 31282 45888 31288
rect 44294 30492 44602 30501
rect 44294 30490 44300 30492
rect 44356 30490 44380 30492
rect 44436 30490 44460 30492
rect 44516 30490 44540 30492
rect 44596 30490 44602 30492
rect 44356 30438 44358 30490
rect 44538 30438 44540 30490
rect 44294 30436 44300 30438
rect 44356 30436 44380 30438
rect 44436 30436 44460 30438
rect 44516 30436 44540 30438
rect 44596 30436 44602 30438
rect 44294 30427 44602 30436
rect 44294 29404 44602 29413
rect 44294 29402 44300 29404
rect 44356 29402 44380 29404
rect 44436 29402 44460 29404
rect 44516 29402 44540 29404
rect 44596 29402 44602 29404
rect 44356 29350 44358 29402
rect 44538 29350 44540 29402
rect 44294 29348 44300 29350
rect 44356 29348 44380 29350
rect 44436 29348 44460 29350
rect 44516 29348 44540 29350
rect 44596 29348 44602 29350
rect 44294 29339 44602 29348
rect 44294 28316 44602 28325
rect 44294 28314 44300 28316
rect 44356 28314 44380 28316
rect 44436 28314 44460 28316
rect 44516 28314 44540 28316
rect 44596 28314 44602 28316
rect 44356 28262 44358 28314
rect 44538 28262 44540 28314
rect 44294 28260 44300 28262
rect 44356 28260 44380 28262
rect 44436 28260 44460 28262
rect 44516 28260 44540 28262
rect 44596 28260 44602 28262
rect 44294 28251 44602 28260
rect 45848 27402 45876 31282
rect 51518 31036 51826 31045
rect 51518 31034 51524 31036
rect 51580 31034 51604 31036
rect 51660 31034 51684 31036
rect 51740 31034 51764 31036
rect 51820 31034 51826 31036
rect 51580 30982 51582 31034
rect 51762 30982 51764 31034
rect 51518 30980 51524 30982
rect 51580 30980 51604 30982
rect 51660 30980 51684 30982
rect 51740 30980 51764 30982
rect 51820 30980 51826 30982
rect 51518 30971 51826 30980
rect 51518 29948 51826 29957
rect 51518 29946 51524 29948
rect 51580 29946 51604 29948
rect 51660 29946 51684 29948
rect 51740 29946 51764 29948
rect 51820 29946 51826 29948
rect 51580 29894 51582 29946
rect 51762 29894 51764 29946
rect 51518 29892 51524 29894
rect 51580 29892 51604 29894
rect 51660 29892 51684 29894
rect 51740 29892 51764 29894
rect 51820 29892 51826 29894
rect 51518 29883 51826 29892
rect 51518 28860 51826 28869
rect 51518 28858 51524 28860
rect 51580 28858 51604 28860
rect 51660 28858 51684 28860
rect 51740 28858 51764 28860
rect 51820 28858 51826 28860
rect 51580 28806 51582 28858
rect 51762 28806 51764 28858
rect 51518 28804 51524 28806
rect 51580 28804 51604 28806
rect 51660 28804 51684 28806
rect 51740 28804 51764 28806
rect 51820 28804 51826 28806
rect 51518 28795 51826 28804
rect 51518 27772 51826 27781
rect 51518 27770 51524 27772
rect 51580 27770 51604 27772
rect 51660 27770 51684 27772
rect 51740 27770 51764 27772
rect 51820 27770 51826 27772
rect 51580 27718 51582 27770
rect 51762 27718 51764 27770
rect 51518 27716 51524 27718
rect 51580 27716 51604 27718
rect 51660 27716 51684 27718
rect 51740 27716 51764 27718
rect 51820 27716 51826 27718
rect 51518 27707 51826 27716
rect 45836 27396 45888 27402
rect 45836 27338 45888 27344
rect 44294 27228 44602 27237
rect 44294 27226 44300 27228
rect 44356 27226 44380 27228
rect 44436 27226 44460 27228
rect 44516 27226 44540 27228
rect 44596 27226 44602 27228
rect 44356 27174 44358 27226
rect 44538 27174 44540 27226
rect 44294 27172 44300 27174
rect 44356 27172 44380 27174
rect 44436 27172 44460 27174
rect 44516 27172 44540 27174
rect 44596 27172 44602 27174
rect 44294 27163 44602 27172
rect 51518 26684 51826 26693
rect 51518 26682 51524 26684
rect 51580 26682 51604 26684
rect 51660 26682 51684 26684
rect 51740 26682 51764 26684
rect 51820 26682 51826 26684
rect 51580 26630 51582 26682
rect 51762 26630 51764 26682
rect 51518 26628 51524 26630
rect 51580 26628 51604 26630
rect 51660 26628 51684 26630
rect 51740 26628 51764 26630
rect 51820 26628 51826 26630
rect 51518 26619 51826 26628
rect 44294 26140 44602 26149
rect 44294 26138 44300 26140
rect 44356 26138 44380 26140
rect 44436 26138 44460 26140
rect 44516 26138 44540 26140
rect 44596 26138 44602 26140
rect 44356 26086 44358 26138
rect 44538 26086 44540 26138
rect 44294 26084 44300 26086
rect 44356 26084 44380 26086
rect 44436 26084 44460 26086
rect 44516 26084 44540 26086
rect 44596 26084 44602 26086
rect 44294 26075 44602 26084
rect 51518 25596 51826 25605
rect 51518 25594 51524 25596
rect 51580 25594 51604 25596
rect 51660 25594 51684 25596
rect 51740 25594 51764 25596
rect 51820 25594 51826 25596
rect 51580 25542 51582 25594
rect 51762 25542 51764 25594
rect 51518 25540 51524 25542
rect 51580 25540 51604 25542
rect 51660 25540 51684 25542
rect 51740 25540 51764 25542
rect 51820 25540 51826 25542
rect 51518 25531 51826 25540
rect 44294 25052 44602 25061
rect 44294 25050 44300 25052
rect 44356 25050 44380 25052
rect 44436 25050 44460 25052
rect 44516 25050 44540 25052
rect 44596 25050 44602 25052
rect 44356 24998 44358 25050
rect 44538 24998 44540 25050
rect 44294 24996 44300 24998
rect 44356 24996 44380 24998
rect 44436 24996 44460 24998
rect 44516 24996 44540 24998
rect 44596 24996 44602 24998
rect 44294 24987 44602 24996
rect 51518 24508 51826 24517
rect 51518 24506 51524 24508
rect 51580 24506 51604 24508
rect 51660 24506 51684 24508
rect 51740 24506 51764 24508
rect 51820 24506 51826 24508
rect 51580 24454 51582 24506
rect 51762 24454 51764 24506
rect 51518 24452 51524 24454
rect 51580 24452 51604 24454
rect 51660 24452 51684 24454
rect 51740 24452 51764 24454
rect 51820 24452 51826 24454
rect 51518 24443 51826 24452
rect 48320 24132 48372 24138
rect 48320 24074 48372 24080
rect 47584 24064 47636 24070
rect 47584 24006 47636 24012
rect 44294 23964 44602 23973
rect 44294 23962 44300 23964
rect 44356 23962 44380 23964
rect 44436 23962 44460 23964
rect 44516 23962 44540 23964
rect 44596 23962 44602 23964
rect 44356 23910 44358 23962
rect 44538 23910 44540 23962
rect 44294 23908 44300 23910
rect 44356 23908 44380 23910
rect 44436 23908 44460 23910
rect 44516 23908 44540 23910
rect 44596 23908 44602 23910
rect 44294 23899 44602 23908
rect 47596 23866 47624 24006
rect 47584 23860 47636 23866
rect 47584 23802 47636 23808
rect 47492 23656 47544 23662
rect 47492 23598 47544 23604
rect 46572 22976 46624 22982
rect 46572 22918 46624 22924
rect 47400 22976 47452 22982
rect 47400 22918 47452 22924
rect 44294 22876 44602 22885
rect 44294 22874 44300 22876
rect 44356 22874 44380 22876
rect 44436 22874 44460 22876
rect 44516 22874 44540 22876
rect 44596 22874 44602 22876
rect 44356 22822 44358 22874
rect 44538 22822 44540 22874
rect 44294 22820 44300 22822
rect 44356 22820 44380 22822
rect 44436 22820 44460 22822
rect 44516 22820 44540 22822
rect 44596 22820 44602 22822
rect 44294 22811 44602 22820
rect 45652 22704 45704 22710
rect 45652 22646 45704 22652
rect 45284 22568 45336 22574
rect 45284 22510 45336 22516
rect 44916 22160 44968 22166
rect 44916 22102 44968 22108
rect 44088 22024 44140 22030
rect 44088 21966 44140 21972
rect 43996 21072 44048 21078
rect 43996 21014 44048 21020
rect 44008 20466 44036 21014
rect 44100 20874 44128 21966
rect 44180 21888 44232 21894
rect 44180 21830 44232 21836
rect 44192 20942 44220 21830
rect 44294 21788 44602 21797
rect 44294 21786 44300 21788
rect 44356 21786 44380 21788
rect 44436 21786 44460 21788
rect 44516 21786 44540 21788
rect 44596 21786 44602 21788
rect 44356 21734 44358 21786
rect 44538 21734 44540 21786
rect 44294 21732 44300 21734
rect 44356 21732 44380 21734
rect 44436 21732 44460 21734
rect 44516 21732 44540 21734
rect 44596 21732 44602 21734
rect 44294 21723 44602 21732
rect 44272 21072 44324 21078
rect 44272 21014 44324 21020
rect 44824 21072 44876 21078
rect 44824 21014 44876 21020
rect 44180 20936 44232 20942
rect 44180 20878 44232 20884
rect 44088 20868 44140 20874
rect 44088 20810 44140 20816
rect 43996 20460 44048 20466
rect 43996 20402 44048 20408
rect 44008 19378 44036 20402
rect 43996 19372 44048 19378
rect 43996 19314 44048 19320
rect 44008 18766 44036 19314
rect 44192 18766 44220 20878
rect 44284 20806 44312 21014
rect 44732 20868 44784 20874
rect 44732 20810 44784 20816
rect 44272 20800 44324 20806
rect 44272 20742 44324 20748
rect 44640 20800 44692 20806
rect 44640 20742 44692 20748
rect 44294 20700 44602 20709
rect 44294 20698 44300 20700
rect 44356 20698 44380 20700
rect 44436 20698 44460 20700
rect 44516 20698 44540 20700
rect 44596 20698 44602 20700
rect 44356 20646 44358 20698
rect 44538 20646 44540 20698
rect 44294 20644 44300 20646
rect 44356 20644 44380 20646
rect 44436 20644 44460 20646
rect 44516 20644 44540 20646
rect 44596 20644 44602 20646
rect 44294 20635 44602 20644
rect 44652 20466 44680 20742
rect 44640 20460 44692 20466
rect 44640 20402 44692 20408
rect 44652 19854 44680 20402
rect 44744 20262 44772 20810
rect 44732 20256 44784 20262
rect 44732 20198 44784 20204
rect 44640 19848 44692 19854
rect 44640 19790 44692 19796
rect 44294 19612 44602 19621
rect 44294 19610 44300 19612
rect 44356 19610 44380 19612
rect 44436 19610 44460 19612
rect 44516 19610 44540 19612
rect 44596 19610 44602 19612
rect 44356 19558 44358 19610
rect 44538 19558 44540 19610
rect 44294 19556 44300 19558
rect 44356 19556 44380 19558
rect 44436 19556 44460 19558
rect 44516 19556 44540 19558
rect 44596 19556 44602 19558
rect 44294 19547 44602 19556
rect 44652 19378 44680 19790
rect 44744 19718 44772 20198
rect 44732 19712 44784 19718
rect 44732 19654 44784 19660
rect 44640 19372 44692 19378
rect 44640 19314 44692 19320
rect 44640 19168 44692 19174
rect 44744 19156 44772 19654
rect 44692 19128 44772 19156
rect 44640 19110 44692 19116
rect 43996 18760 44048 18766
rect 43996 18702 44048 18708
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 44652 18698 44680 19110
rect 44640 18692 44692 18698
rect 44640 18634 44692 18640
rect 44294 18524 44602 18533
rect 44294 18522 44300 18524
rect 44356 18522 44380 18524
rect 44436 18522 44460 18524
rect 44516 18522 44540 18524
rect 44596 18522 44602 18524
rect 44356 18470 44358 18522
rect 44538 18470 44540 18522
rect 44294 18468 44300 18470
rect 44356 18468 44380 18470
rect 44436 18468 44460 18470
rect 44516 18468 44540 18470
rect 44596 18468 44602 18470
rect 44294 18459 44602 18468
rect 44652 18358 44680 18634
rect 44640 18352 44692 18358
rect 44640 18294 44692 18300
rect 43996 18080 44048 18086
rect 43996 18022 44048 18028
rect 43904 16448 43956 16454
rect 43904 16390 43956 16396
rect 44008 14550 44036 18022
rect 44180 17672 44232 17678
rect 44180 17614 44232 17620
rect 44192 17338 44220 17614
rect 44294 17436 44602 17445
rect 44294 17434 44300 17436
rect 44356 17434 44380 17436
rect 44436 17434 44460 17436
rect 44516 17434 44540 17436
rect 44596 17434 44602 17436
rect 44356 17382 44358 17434
rect 44538 17382 44540 17434
rect 44294 17380 44300 17382
rect 44356 17380 44380 17382
rect 44436 17380 44460 17382
rect 44516 17380 44540 17382
rect 44596 17380 44602 17382
rect 44294 17371 44602 17380
rect 44836 17338 44864 21014
rect 44928 20874 44956 22102
rect 45296 22098 45324 22510
rect 45664 22234 45692 22646
rect 46584 22506 46612 22918
rect 46572 22500 46624 22506
rect 46572 22442 46624 22448
rect 45652 22228 45704 22234
rect 45652 22170 45704 22176
rect 45284 22092 45336 22098
rect 45284 22034 45336 22040
rect 45296 21962 45324 22034
rect 45376 22024 45428 22030
rect 45376 21966 45428 21972
rect 45284 21956 45336 21962
rect 45284 21898 45336 21904
rect 45008 21888 45060 21894
rect 45008 21830 45060 21836
rect 45020 21554 45048 21830
rect 45388 21690 45416 21966
rect 45376 21684 45428 21690
rect 45376 21626 45428 21632
rect 45664 21622 45692 22170
rect 46204 22024 46256 22030
rect 46204 21966 46256 21972
rect 45744 21888 45796 21894
rect 45744 21830 45796 21836
rect 45652 21616 45704 21622
rect 45652 21558 45704 21564
rect 45008 21548 45060 21554
rect 45008 21490 45060 21496
rect 44916 20868 44968 20874
rect 44916 20810 44968 20816
rect 45376 20392 45428 20398
rect 45376 20334 45428 20340
rect 45388 19378 45416 20334
rect 45376 19372 45428 19378
rect 45376 19314 45428 19320
rect 45664 18902 45692 21558
rect 45756 20942 45784 21830
rect 46216 21146 46244 21966
rect 46584 21894 46612 22442
rect 46848 22432 46900 22438
rect 46848 22374 46900 22380
rect 46572 21888 46624 21894
rect 46572 21830 46624 21836
rect 46204 21140 46256 21146
rect 46204 21082 46256 21088
rect 46860 21078 46888 22374
rect 47216 22092 47268 22098
rect 47216 22034 47268 22040
rect 47228 21146 47256 22034
rect 47412 21486 47440 22918
rect 47504 21690 47532 23598
rect 47596 23186 47624 23802
rect 47584 23180 47636 23186
rect 47584 23122 47636 23128
rect 47768 23112 47820 23118
rect 47768 23054 47820 23060
rect 47676 22568 47728 22574
rect 47676 22510 47728 22516
rect 47582 21992 47638 22001
rect 47582 21927 47638 21936
rect 47596 21894 47624 21927
rect 47584 21888 47636 21894
rect 47584 21830 47636 21836
rect 47492 21684 47544 21690
rect 47492 21626 47544 21632
rect 47400 21480 47452 21486
rect 47400 21422 47452 21428
rect 47400 21344 47452 21350
rect 47400 21286 47452 21292
rect 47216 21140 47268 21146
rect 47216 21082 47268 21088
rect 46848 21072 46900 21078
rect 46848 21014 46900 21020
rect 47412 20942 47440 21286
rect 47504 21146 47532 21626
rect 47688 21554 47716 22510
rect 47780 22030 47808 23054
rect 48332 22710 48360 24074
rect 48596 23656 48648 23662
rect 48596 23598 48648 23604
rect 48608 23186 48636 23598
rect 51518 23420 51826 23429
rect 51518 23418 51524 23420
rect 51580 23418 51604 23420
rect 51660 23418 51684 23420
rect 51740 23418 51764 23420
rect 51820 23418 51826 23420
rect 51580 23366 51582 23418
rect 51762 23366 51764 23418
rect 51518 23364 51524 23366
rect 51580 23364 51604 23366
rect 51660 23364 51684 23366
rect 51740 23364 51764 23366
rect 51820 23364 51826 23366
rect 51518 23355 51826 23364
rect 48596 23180 48648 23186
rect 48596 23122 48648 23128
rect 48320 22704 48372 22710
rect 48320 22646 48372 22652
rect 48608 22574 48636 23122
rect 51908 22636 51960 22642
rect 51908 22578 51960 22584
rect 48596 22568 48648 22574
rect 48596 22510 48648 22516
rect 49148 22568 49200 22574
rect 49148 22510 49200 22516
rect 48044 22500 48096 22506
rect 48044 22442 48096 22448
rect 47768 22024 47820 22030
rect 47768 21966 47820 21972
rect 47780 21554 47808 21966
rect 47676 21548 47728 21554
rect 47676 21490 47728 21496
rect 47768 21548 47820 21554
rect 47768 21490 47820 21496
rect 47768 21412 47820 21418
rect 47768 21354 47820 21360
rect 47492 21140 47544 21146
rect 47492 21082 47544 21088
rect 47780 20942 47808 21354
rect 45744 20936 45796 20942
rect 45744 20878 45796 20884
rect 47400 20936 47452 20942
rect 47400 20878 47452 20884
rect 47676 20936 47728 20942
rect 47676 20878 47728 20884
rect 47768 20936 47820 20942
rect 47768 20878 47820 20884
rect 45756 20466 45784 20878
rect 46480 20800 46532 20806
rect 46480 20742 46532 20748
rect 45744 20460 45796 20466
rect 45744 20402 45796 20408
rect 46296 20460 46348 20466
rect 46296 20402 46348 20408
rect 45756 19854 45784 20402
rect 45744 19848 45796 19854
rect 45744 19790 45796 19796
rect 45756 19378 45784 19790
rect 46308 19378 46336 20402
rect 46492 19786 46520 20742
rect 47492 20460 47544 20466
rect 47492 20402 47544 20408
rect 46572 20256 46624 20262
rect 46572 20198 46624 20204
rect 46480 19780 46532 19786
rect 46480 19722 46532 19728
rect 45744 19372 45796 19378
rect 45744 19314 45796 19320
rect 46296 19372 46348 19378
rect 46296 19314 46348 19320
rect 45652 18896 45704 18902
rect 45652 18838 45704 18844
rect 46308 18766 46336 19314
rect 46492 19310 46520 19722
rect 46584 19718 46612 20198
rect 46572 19712 46624 19718
rect 46572 19654 46624 19660
rect 46584 19446 46612 19654
rect 46572 19440 46624 19446
rect 46572 19382 46624 19388
rect 46480 19304 46532 19310
rect 46480 19246 46532 19252
rect 46492 19174 46520 19246
rect 46480 19168 46532 19174
rect 46480 19110 46532 19116
rect 46296 18760 46348 18766
rect 46296 18702 46348 18708
rect 45928 18692 45980 18698
rect 45928 18634 45980 18640
rect 45560 18352 45612 18358
rect 45560 18294 45612 18300
rect 45836 18352 45888 18358
rect 45836 18294 45888 18300
rect 45008 17672 45060 17678
rect 45008 17614 45060 17620
rect 44180 17332 44232 17338
rect 44180 17274 44232 17280
rect 44824 17332 44876 17338
rect 44824 17274 44876 17280
rect 44088 16788 44140 16794
rect 44088 16730 44140 16736
rect 44100 16522 44128 16730
rect 44192 16658 44220 17274
rect 44272 16788 44324 16794
rect 44272 16730 44324 16736
rect 44180 16652 44232 16658
rect 44180 16594 44232 16600
rect 44284 16538 44312 16730
rect 44916 16720 44968 16726
rect 44916 16662 44968 16668
rect 44640 16652 44692 16658
rect 44640 16594 44692 16600
rect 44088 16516 44140 16522
rect 44088 16458 44140 16464
rect 44192 16510 44312 16538
rect 44192 16402 44220 16510
rect 44100 16374 44220 16402
rect 44100 15502 44128 16374
rect 44294 16348 44602 16357
rect 44294 16346 44300 16348
rect 44356 16346 44380 16348
rect 44436 16346 44460 16348
rect 44516 16346 44540 16348
rect 44596 16346 44602 16348
rect 44356 16294 44358 16346
rect 44538 16294 44540 16346
rect 44294 16292 44300 16294
rect 44356 16292 44380 16294
rect 44436 16292 44460 16294
rect 44516 16292 44540 16294
rect 44596 16292 44602 16294
rect 44294 16283 44602 16292
rect 44180 16040 44232 16046
rect 44180 15982 44232 15988
rect 44088 15496 44140 15502
rect 44088 15438 44140 15444
rect 44192 14550 44220 15982
rect 44652 15638 44680 16594
rect 44732 15904 44784 15910
rect 44732 15846 44784 15852
rect 44640 15632 44692 15638
rect 44640 15574 44692 15580
rect 44640 15360 44692 15366
rect 44640 15302 44692 15308
rect 44294 15260 44602 15269
rect 44294 15258 44300 15260
rect 44356 15258 44380 15260
rect 44436 15258 44460 15260
rect 44516 15258 44540 15260
rect 44596 15258 44602 15260
rect 44356 15206 44358 15258
rect 44538 15206 44540 15258
rect 44294 15204 44300 15206
rect 44356 15204 44380 15206
rect 44436 15204 44460 15206
rect 44516 15204 44540 15206
rect 44596 15204 44602 15206
rect 44294 15195 44602 15204
rect 44652 14890 44680 15302
rect 44744 15094 44772 15846
rect 44824 15360 44876 15366
rect 44824 15302 44876 15308
rect 44732 15088 44784 15094
rect 44732 15030 44784 15036
rect 44836 14958 44864 15302
rect 44824 14952 44876 14958
rect 44824 14894 44876 14900
rect 44640 14884 44692 14890
rect 44640 14826 44692 14832
rect 43996 14544 44048 14550
rect 43996 14486 44048 14492
rect 44180 14544 44232 14550
rect 44180 14486 44232 14492
rect 44008 14278 44036 14486
rect 44652 14414 44680 14826
rect 44928 14822 44956 16662
rect 45020 15910 45048 17614
rect 45192 17604 45244 17610
rect 45192 17546 45244 17552
rect 45204 17241 45232 17546
rect 45190 17232 45246 17241
rect 45190 17167 45246 17176
rect 45572 16182 45600 18294
rect 45652 17128 45704 17134
rect 45652 17070 45704 17076
rect 45664 16250 45692 17070
rect 45848 16454 45876 18294
rect 45940 18222 45968 18634
rect 45928 18216 45980 18222
rect 45928 18158 45980 18164
rect 45940 17610 45968 18158
rect 45928 17604 45980 17610
rect 45928 17546 45980 17552
rect 45940 17134 45968 17546
rect 45928 17128 45980 17134
rect 45928 17070 45980 17076
rect 45836 16448 45888 16454
rect 45836 16390 45888 16396
rect 45652 16244 45704 16250
rect 45652 16186 45704 16192
rect 45192 16176 45244 16182
rect 45192 16118 45244 16124
rect 45560 16176 45612 16182
rect 45560 16118 45612 16124
rect 45008 15904 45060 15910
rect 45008 15846 45060 15852
rect 45008 15496 45060 15502
rect 45008 15438 45060 15444
rect 45020 15162 45048 15438
rect 45008 15156 45060 15162
rect 45008 15098 45060 15104
rect 45100 14952 45152 14958
rect 45100 14894 45152 14900
rect 44916 14816 44968 14822
rect 44916 14758 44968 14764
rect 44928 14482 44956 14758
rect 45112 14618 45140 14894
rect 45100 14612 45152 14618
rect 45100 14554 45152 14560
rect 44916 14476 44968 14482
rect 44916 14418 44968 14424
rect 44640 14408 44692 14414
rect 44640 14350 44692 14356
rect 44824 14340 44876 14346
rect 44824 14282 44876 14288
rect 43996 14272 44048 14278
rect 43996 14214 44048 14220
rect 44008 14074 44036 14214
rect 44294 14172 44602 14181
rect 44294 14170 44300 14172
rect 44356 14170 44380 14172
rect 44436 14170 44460 14172
rect 44516 14170 44540 14172
rect 44596 14170 44602 14172
rect 44356 14118 44358 14170
rect 44538 14118 44540 14170
rect 44294 14116 44300 14118
rect 44356 14116 44380 14118
rect 44436 14116 44460 14118
rect 44516 14116 44540 14118
rect 44596 14116 44602 14118
rect 44294 14107 44602 14116
rect 43996 14068 44048 14074
rect 43996 14010 44048 14016
rect 44008 13530 44036 14010
rect 44836 14006 44864 14282
rect 44928 14006 44956 14418
rect 45204 14346 45232 16118
rect 45848 16114 45876 16390
rect 45836 16108 45888 16114
rect 45836 16050 45888 16056
rect 45560 15904 45612 15910
rect 45560 15846 45612 15852
rect 45468 15156 45520 15162
rect 45468 15098 45520 15104
rect 45376 14544 45428 14550
rect 45376 14486 45428 14492
rect 45192 14340 45244 14346
rect 45192 14282 45244 14288
rect 44824 14000 44876 14006
rect 44824 13942 44876 13948
rect 44916 14000 44968 14006
rect 44916 13942 44968 13948
rect 45100 14000 45152 14006
rect 45100 13942 45152 13948
rect 43996 13524 44048 13530
rect 43996 13466 44048 13472
rect 44836 13326 44864 13942
rect 44824 13320 44876 13326
rect 44824 13262 44876 13268
rect 44916 13184 44968 13190
rect 44916 13126 44968 13132
rect 44294 13084 44602 13093
rect 44294 13082 44300 13084
rect 44356 13082 44380 13084
rect 44436 13082 44460 13084
rect 44516 13082 44540 13084
rect 44596 13082 44602 13084
rect 44356 13030 44358 13082
rect 44538 13030 44540 13082
rect 44294 13028 44300 13030
rect 44356 13028 44380 13030
rect 44436 13028 44460 13030
rect 44516 13028 44540 13030
rect 44596 13028 44602 13030
rect 44294 13019 44602 13028
rect 44928 12850 44956 13126
rect 44732 12844 44784 12850
rect 44732 12786 44784 12792
rect 44916 12844 44968 12850
rect 44916 12786 44968 12792
rect 44744 12434 44772 12786
rect 45112 12434 45140 13942
rect 45192 13932 45244 13938
rect 45192 13874 45244 13880
rect 45204 13394 45232 13874
rect 45192 13388 45244 13394
rect 45192 13330 45244 13336
rect 45204 12968 45232 13330
rect 45388 13274 45416 14486
rect 45480 14074 45508 15098
rect 45572 14414 45600 15846
rect 45940 15570 45968 17070
rect 46492 16114 46520 19110
rect 47400 18692 47452 18698
rect 47400 18634 47452 18640
rect 46846 18320 46902 18329
rect 46846 18255 46902 18264
rect 46860 18222 46888 18255
rect 46848 18216 46900 18222
rect 46848 18158 46900 18164
rect 47032 18216 47084 18222
rect 47032 18158 47084 18164
rect 46756 18148 46808 18154
rect 46756 18090 46808 18096
rect 46768 17338 46796 18090
rect 46756 17332 46808 17338
rect 46756 17274 46808 17280
rect 47044 16794 47072 18158
rect 47412 17746 47440 18634
rect 47400 17740 47452 17746
rect 47400 17682 47452 17688
rect 47032 16788 47084 16794
rect 47032 16730 47084 16736
rect 46848 16244 46900 16250
rect 46848 16186 46900 16192
rect 46480 16108 46532 16114
rect 46480 16050 46532 16056
rect 46020 15972 46072 15978
rect 46020 15914 46072 15920
rect 46032 15570 46060 15914
rect 45928 15564 45980 15570
rect 45928 15506 45980 15512
rect 46020 15564 46072 15570
rect 46020 15506 46072 15512
rect 45940 15366 45968 15506
rect 45928 15360 45980 15366
rect 45928 15302 45980 15308
rect 45836 14952 45888 14958
rect 45836 14894 45888 14900
rect 45848 14550 45876 14894
rect 45836 14544 45888 14550
rect 45836 14486 45888 14492
rect 45560 14408 45612 14414
rect 45560 14350 45612 14356
rect 45836 14340 45888 14346
rect 45836 14282 45888 14288
rect 45468 14068 45520 14074
rect 45468 14010 45520 14016
rect 45480 13530 45508 14010
rect 45848 13938 45876 14282
rect 45928 14272 45980 14278
rect 45928 14214 45980 14220
rect 45836 13932 45888 13938
rect 45836 13874 45888 13880
rect 45940 13802 45968 14214
rect 46032 13938 46060 15506
rect 46112 15428 46164 15434
rect 46112 15370 46164 15376
rect 46124 14618 46152 15370
rect 46112 14612 46164 14618
rect 46112 14554 46164 14560
rect 46204 14476 46256 14482
rect 46204 14418 46256 14424
rect 46296 14476 46348 14482
rect 46296 14418 46348 14424
rect 46020 13932 46072 13938
rect 46020 13874 46072 13880
rect 46216 13870 46244 14418
rect 46308 14074 46336 14418
rect 46296 14068 46348 14074
rect 46296 14010 46348 14016
rect 46204 13864 46256 13870
rect 46204 13806 46256 13812
rect 45928 13796 45980 13802
rect 45928 13738 45980 13744
rect 45468 13524 45520 13530
rect 45468 13466 45520 13472
rect 45560 13320 45612 13326
rect 45480 13280 45560 13308
rect 45480 13274 45508 13280
rect 45388 13258 45508 13274
rect 45560 13262 45612 13268
rect 46296 13320 46348 13326
rect 46296 13262 46348 13268
rect 45376 13252 45508 13258
rect 45428 13246 45508 13252
rect 45376 13194 45428 13200
rect 45204 12940 45324 12968
rect 45192 12844 45244 12850
rect 45192 12786 45244 12792
rect 44744 12406 44864 12434
rect 43628 12164 43680 12170
rect 43628 12106 43680 12112
rect 43640 11744 43668 12106
rect 44180 12096 44232 12102
rect 44180 12038 44232 12044
rect 44192 11830 44220 12038
rect 44294 11996 44602 12005
rect 44294 11994 44300 11996
rect 44356 11994 44380 11996
rect 44436 11994 44460 11996
rect 44516 11994 44540 11996
rect 44596 11994 44602 11996
rect 44356 11942 44358 11994
rect 44538 11942 44540 11994
rect 44294 11940 44300 11942
rect 44356 11940 44380 11942
rect 44436 11940 44460 11942
rect 44516 11940 44540 11942
rect 44596 11940 44602 11942
rect 44294 11931 44602 11940
rect 43812 11824 43864 11830
rect 43812 11766 43864 11772
rect 44180 11824 44232 11830
rect 44180 11766 44232 11772
rect 43720 11756 43772 11762
rect 43640 11716 43720 11744
rect 43720 11698 43772 11704
rect 43444 11688 43496 11694
rect 43444 11630 43496 11636
rect 42708 11348 42760 11354
rect 42708 11290 42760 11296
rect 42524 10668 42576 10674
rect 42524 10610 42576 10616
rect 42616 10668 42668 10674
rect 42616 10610 42668 10616
rect 42536 9994 42564 10610
rect 42524 9988 42576 9994
rect 42524 9930 42576 9936
rect 42340 9036 42392 9042
rect 42340 8978 42392 8984
rect 42352 7954 42380 8978
rect 42536 8922 42564 9930
rect 42628 9722 42656 10610
rect 42720 9994 42748 11290
rect 43456 10810 43484 11630
rect 43824 11286 43852 11766
rect 43812 11280 43864 11286
rect 43812 11222 43864 11228
rect 43536 11008 43588 11014
rect 43536 10950 43588 10956
rect 43444 10804 43496 10810
rect 43444 10746 43496 10752
rect 43548 10674 43576 10950
rect 43824 10674 43852 11222
rect 44294 10908 44602 10917
rect 44294 10906 44300 10908
rect 44356 10906 44380 10908
rect 44436 10906 44460 10908
rect 44516 10906 44540 10908
rect 44596 10906 44602 10908
rect 44356 10854 44358 10906
rect 44538 10854 44540 10906
rect 44294 10852 44300 10854
rect 44356 10852 44380 10854
rect 44436 10852 44460 10854
rect 44516 10852 44540 10854
rect 44596 10852 44602 10854
rect 44294 10843 44602 10852
rect 43536 10668 43588 10674
rect 43536 10610 43588 10616
rect 43812 10668 43864 10674
rect 43812 10610 43864 10616
rect 43548 10470 43576 10610
rect 43536 10464 43588 10470
rect 43536 10406 43588 10412
rect 42708 9988 42760 9994
rect 42708 9930 42760 9936
rect 43548 9722 43576 10406
rect 44180 9920 44232 9926
rect 44180 9862 44232 9868
rect 42616 9716 42668 9722
rect 42616 9658 42668 9664
rect 43536 9716 43588 9722
rect 43536 9658 43588 9664
rect 42444 8906 42564 8922
rect 42432 8900 42564 8906
rect 42484 8894 42564 8900
rect 42432 8842 42484 8848
rect 42628 8430 42656 9658
rect 42892 9376 42944 9382
rect 42892 9318 42944 9324
rect 42904 9178 42932 9318
rect 42892 9172 42944 9178
rect 42892 9114 42944 9120
rect 44192 9058 44220 9862
rect 44294 9820 44602 9829
rect 44294 9818 44300 9820
rect 44356 9818 44380 9820
rect 44436 9818 44460 9820
rect 44516 9818 44540 9820
rect 44596 9818 44602 9820
rect 44356 9766 44358 9818
rect 44538 9766 44540 9818
rect 44294 9764 44300 9766
rect 44356 9764 44380 9766
rect 44436 9764 44460 9766
rect 44516 9764 44540 9766
rect 44596 9764 44602 9766
rect 44294 9755 44602 9764
rect 44836 9654 44864 12406
rect 44928 12406 45140 12434
rect 44928 11150 44956 12406
rect 45204 11830 45232 12786
rect 45296 12782 45324 12940
rect 45284 12776 45336 12782
rect 45284 12718 45336 12724
rect 45284 12640 45336 12646
rect 45284 12582 45336 12588
rect 45192 11824 45244 11830
rect 45192 11766 45244 11772
rect 45100 11688 45152 11694
rect 45100 11630 45152 11636
rect 45112 11354 45140 11630
rect 45100 11348 45152 11354
rect 45100 11290 45152 11296
rect 45296 11218 45324 12582
rect 46308 12442 46336 13262
rect 46492 12646 46520 16050
rect 46756 16040 46808 16046
rect 46756 15982 46808 15988
rect 46664 14408 46716 14414
rect 46664 14350 46716 14356
rect 46676 14074 46704 14350
rect 46664 14068 46716 14074
rect 46664 14010 46716 14016
rect 46768 12850 46796 15982
rect 46860 15094 46888 16186
rect 47504 15434 47532 20402
rect 47688 19310 47716 20878
rect 47780 20466 47808 20878
rect 47768 20460 47820 20466
rect 47768 20402 47820 20408
rect 47952 19372 48004 19378
rect 47952 19314 48004 19320
rect 47676 19304 47728 19310
rect 47676 19246 47728 19252
rect 47676 18760 47728 18766
rect 47676 18702 47728 18708
rect 47688 17746 47716 18702
rect 47676 17740 47728 17746
rect 47676 17682 47728 17688
rect 47768 17196 47820 17202
rect 47768 17138 47820 17144
rect 47676 16992 47728 16998
rect 47676 16934 47728 16940
rect 47688 15706 47716 16934
rect 47780 16658 47808 17138
rect 47768 16652 47820 16658
rect 47768 16594 47820 16600
rect 47676 15700 47728 15706
rect 47676 15642 47728 15648
rect 46940 15428 46992 15434
rect 46940 15370 46992 15376
rect 47492 15428 47544 15434
rect 47492 15370 47544 15376
rect 46848 15088 46900 15094
rect 46848 15030 46900 15036
rect 46860 14414 46888 15030
rect 46848 14408 46900 14414
rect 46848 14350 46900 14356
rect 46756 12844 46808 12850
rect 46756 12786 46808 12792
rect 46952 12714 46980 15370
rect 47308 15360 47360 15366
rect 47308 15302 47360 15308
rect 47216 14272 47268 14278
rect 47216 14214 47268 14220
rect 47228 14006 47256 14214
rect 47216 14000 47268 14006
rect 47216 13942 47268 13948
rect 47216 13320 47268 13326
rect 47320 13308 47348 15302
rect 47492 15020 47544 15026
rect 47492 14962 47544 14968
rect 47504 14278 47532 14962
rect 47492 14272 47544 14278
rect 47492 14214 47544 14220
rect 47504 13326 47532 14214
rect 47268 13280 47348 13308
rect 47492 13320 47544 13326
rect 47216 13262 47268 13268
rect 47492 13262 47544 13268
rect 47032 13184 47084 13190
rect 47032 13126 47084 13132
rect 46940 12708 46992 12714
rect 46940 12650 46992 12656
rect 46480 12640 46532 12646
rect 46480 12582 46532 12588
rect 46296 12436 46348 12442
rect 46296 12378 46348 12384
rect 45376 12164 45428 12170
rect 45376 12106 45428 12112
rect 45388 11898 45416 12106
rect 45376 11892 45428 11898
rect 45376 11834 45428 11840
rect 45376 11552 45428 11558
rect 45376 11494 45428 11500
rect 45468 11552 45520 11558
rect 45468 11494 45520 11500
rect 45388 11354 45416 11494
rect 45376 11348 45428 11354
rect 45376 11290 45428 11296
rect 45284 11212 45336 11218
rect 45284 11154 45336 11160
rect 45480 11150 45508 11494
rect 44916 11144 44968 11150
rect 44916 11086 44968 11092
rect 45468 11144 45520 11150
rect 45468 11086 45520 11092
rect 45376 10464 45428 10470
rect 45376 10406 45428 10412
rect 45560 10464 45612 10470
rect 45560 10406 45612 10412
rect 44824 9648 44876 9654
rect 44824 9590 44876 9596
rect 44732 9580 44784 9586
rect 44732 9522 44784 9528
rect 44100 9030 44220 9058
rect 44100 8974 44128 9030
rect 44088 8968 44140 8974
rect 44088 8910 44140 8916
rect 42892 8832 42944 8838
rect 42892 8774 42944 8780
rect 42904 8634 42932 8774
rect 42892 8628 42944 8634
rect 42892 8570 42944 8576
rect 44100 8514 44128 8910
rect 44180 8900 44232 8906
rect 44180 8842 44232 8848
rect 44192 8616 44220 8842
rect 44294 8732 44602 8741
rect 44294 8730 44300 8732
rect 44356 8730 44380 8732
rect 44436 8730 44460 8732
rect 44516 8730 44540 8732
rect 44596 8730 44602 8732
rect 44356 8678 44358 8730
rect 44538 8678 44540 8730
rect 44294 8676 44300 8678
rect 44356 8676 44380 8678
rect 44436 8676 44460 8678
rect 44516 8676 44540 8678
rect 44596 8676 44602 8678
rect 44294 8667 44602 8676
rect 44744 8634 44772 9522
rect 44732 8628 44784 8634
rect 44192 8588 44404 8616
rect 44100 8486 44220 8514
rect 44376 8498 44404 8588
rect 44732 8570 44784 8576
rect 42616 8424 42668 8430
rect 42616 8366 42668 8372
rect 43076 8288 43128 8294
rect 43074 8256 43076 8265
rect 44192 8276 44220 8486
rect 44364 8492 44416 8498
rect 44364 8434 44416 8440
rect 44640 8492 44692 8498
rect 44640 8434 44692 8440
rect 44272 8288 44324 8294
rect 43128 8256 43130 8265
rect 43074 8191 43130 8200
rect 44192 8248 44272 8276
rect 42340 7948 42392 7954
rect 42340 7890 42392 7896
rect 42352 7410 42380 7890
rect 43168 7812 43220 7818
rect 43168 7754 43220 7760
rect 43180 7478 43208 7754
rect 43168 7472 43220 7478
rect 43168 7414 43220 7420
rect 42340 7404 42392 7410
rect 42340 7346 42392 7352
rect 44088 6792 44140 6798
rect 44088 6734 44140 6740
rect 43076 6724 43128 6730
rect 43076 6666 43128 6672
rect 42892 6656 42944 6662
rect 42892 6598 42944 6604
rect 42984 6656 43036 6662
rect 42984 6598 43036 6604
rect 42904 6322 42932 6598
rect 42996 6322 43024 6598
rect 42892 6316 42944 6322
rect 42892 6258 42944 6264
rect 42984 6316 43036 6322
rect 42984 6258 43036 6264
rect 42904 5642 42932 6258
rect 42996 5846 43024 6258
rect 43088 6118 43116 6666
rect 43996 6316 44048 6322
rect 43996 6258 44048 6264
rect 43628 6180 43680 6186
rect 43628 6122 43680 6128
rect 43076 6112 43128 6118
rect 43076 6054 43128 6060
rect 43536 6112 43588 6118
rect 43536 6054 43588 6060
rect 42984 5840 43036 5846
rect 42984 5782 43036 5788
rect 43548 5642 43576 6054
rect 42892 5636 42944 5642
rect 42892 5578 42944 5584
rect 43444 5636 43496 5642
rect 43444 5578 43496 5584
rect 43536 5636 43588 5642
rect 43536 5578 43588 5584
rect 42708 5568 42760 5574
rect 42708 5510 42760 5516
rect 42432 4684 42484 4690
rect 42432 4626 42484 4632
rect 42062 4584 42118 4593
rect 42062 4519 42118 4528
rect 42444 4146 42472 4626
rect 42432 4140 42484 4146
rect 42432 4082 42484 4088
rect 42720 4078 42748 5510
rect 43076 5228 43128 5234
rect 43076 5170 43128 5176
rect 43088 4078 43116 5170
rect 43456 5166 43484 5578
rect 43444 5160 43496 5166
rect 43444 5102 43496 5108
rect 43548 5030 43576 5578
rect 43536 5024 43588 5030
rect 43536 4966 43588 4972
rect 43640 4554 43668 6122
rect 44008 5574 44036 6258
rect 44100 5710 44128 6734
rect 44088 5704 44140 5710
rect 44088 5646 44140 5652
rect 43996 5568 44048 5574
rect 43996 5510 44048 5516
rect 43628 4548 43680 4554
rect 43628 4490 43680 4496
rect 42708 4072 42760 4078
rect 42708 4014 42760 4020
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 41788 3664 41840 3670
rect 41788 3606 41840 3612
rect 44192 3194 44220 8248
rect 44272 8230 44324 8236
rect 44376 8090 44404 8434
rect 44364 8084 44416 8090
rect 44364 8026 44416 8032
rect 44294 7644 44602 7653
rect 44294 7642 44300 7644
rect 44356 7642 44380 7644
rect 44436 7642 44460 7644
rect 44516 7642 44540 7644
rect 44596 7642 44602 7644
rect 44356 7590 44358 7642
rect 44538 7590 44540 7642
rect 44294 7588 44300 7590
rect 44356 7588 44380 7590
rect 44436 7588 44460 7590
rect 44516 7588 44540 7590
rect 44596 7588 44602 7590
rect 44294 7579 44602 7588
rect 44652 7546 44680 8434
rect 44744 7546 44772 8570
rect 44836 8401 44864 9590
rect 45100 8968 45152 8974
rect 45100 8910 45152 8916
rect 45112 8634 45140 8910
rect 45388 8838 45416 10406
rect 45572 10266 45600 10406
rect 45560 10260 45612 10266
rect 45560 10202 45612 10208
rect 45468 9988 45520 9994
rect 45468 9930 45520 9936
rect 45480 9586 45508 9930
rect 45468 9580 45520 9586
rect 45468 9522 45520 9528
rect 46952 9450 46980 12650
rect 47044 12306 47072 13126
rect 47032 12300 47084 12306
rect 47032 12242 47084 12248
rect 47400 11144 47452 11150
rect 47400 11086 47452 11092
rect 47412 11014 47440 11086
rect 47400 11008 47452 11014
rect 47400 10950 47452 10956
rect 46940 9444 46992 9450
rect 46940 9386 46992 9392
rect 45560 9104 45612 9110
rect 45560 9046 45612 9052
rect 45192 8832 45244 8838
rect 45192 8774 45244 8780
rect 45376 8832 45428 8838
rect 45376 8774 45428 8780
rect 45100 8628 45152 8634
rect 45100 8570 45152 8576
rect 45112 8498 45140 8570
rect 45100 8492 45152 8498
rect 45100 8434 45152 8440
rect 44822 8392 44878 8401
rect 44822 8327 44878 8336
rect 44640 7540 44692 7546
rect 44640 7482 44692 7488
rect 44732 7540 44784 7546
rect 44732 7482 44784 7488
rect 44744 6730 44772 7482
rect 45100 7404 45152 7410
rect 45100 7346 45152 7352
rect 45112 7002 45140 7346
rect 45204 7342 45232 8774
rect 45388 8616 45416 8774
rect 45572 8634 45600 9046
rect 46204 9036 46256 9042
rect 46204 8978 46256 8984
rect 45928 8900 45980 8906
rect 45928 8842 45980 8848
rect 45560 8628 45612 8634
rect 45388 8588 45508 8616
rect 45376 8492 45428 8498
rect 45376 8434 45428 8440
rect 45388 7886 45416 8434
rect 45376 7880 45428 7886
rect 45376 7822 45428 7828
rect 45480 7410 45508 8588
rect 45560 8570 45612 8576
rect 45572 7478 45600 8570
rect 45560 7472 45612 7478
rect 45560 7414 45612 7420
rect 45468 7404 45520 7410
rect 45468 7346 45520 7352
rect 45192 7336 45244 7342
rect 45192 7278 45244 7284
rect 45100 6996 45152 7002
rect 45100 6938 45152 6944
rect 45572 6798 45600 7414
rect 45940 7410 45968 8842
rect 46216 8634 46244 8978
rect 47688 8838 47716 15642
rect 47964 11744 47992 19314
rect 48056 19310 48084 22442
rect 49160 22234 49188 22510
rect 51518 22332 51826 22341
rect 51518 22330 51524 22332
rect 51580 22330 51604 22332
rect 51660 22330 51684 22332
rect 51740 22330 51764 22332
rect 51820 22330 51826 22332
rect 51580 22278 51582 22330
rect 51762 22278 51764 22330
rect 51518 22276 51524 22278
rect 51580 22276 51604 22278
rect 51660 22276 51684 22278
rect 51740 22276 51764 22278
rect 51820 22276 51826 22278
rect 51518 22267 51826 22276
rect 49148 22228 49200 22234
rect 49148 22170 49200 22176
rect 49608 22228 49660 22234
rect 49608 22170 49660 22176
rect 48320 22092 48372 22098
rect 48320 22034 48372 22040
rect 48332 19514 48360 22034
rect 48412 21956 48464 21962
rect 48412 21898 48464 21904
rect 48424 21554 48452 21898
rect 48596 21888 48648 21894
rect 48596 21830 48648 21836
rect 48608 21622 48636 21830
rect 49160 21622 49188 22170
rect 49240 21888 49292 21894
rect 49240 21830 49292 21836
rect 48596 21616 48648 21622
rect 48596 21558 48648 21564
rect 49148 21616 49200 21622
rect 49148 21558 49200 21564
rect 48412 21548 48464 21554
rect 48412 21490 48464 21496
rect 49056 21344 49108 21350
rect 49056 21286 49108 21292
rect 48412 20936 48464 20942
rect 48412 20878 48464 20884
rect 48424 20330 48452 20878
rect 49068 20874 49096 21286
rect 49252 21010 49280 21830
rect 49620 21690 49648 22170
rect 50620 22092 50672 22098
rect 50620 22034 50672 22040
rect 50160 22024 50212 22030
rect 50160 21966 50212 21972
rect 49976 21888 50028 21894
rect 49976 21830 50028 21836
rect 49516 21684 49568 21690
rect 49516 21626 49568 21632
rect 49608 21684 49660 21690
rect 49608 21626 49660 21632
rect 49332 21480 49384 21486
rect 49332 21422 49384 21428
rect 49344 21146 49372 21422
rect 49332 21140 49384 21146
rect 49332 21082 49384 21088
rect 49240 21004 49292 21010
rect 49240 20946 49292 20952
rect 49056 20868 49108 20874
rect 49056 20810 49108 20816
rect 48872 20800 48924 20806
rect 48872 20742 48924 20748
rect 48412 20324 48464 20330
rect 48412 20266 48464 20272
rect 48688 20256 48740 20262
rect 48688 20198 48740 20204
rect 48320 19508 48372 19514
rect 48320 19450 48372 19456
rect 48044 19304 48096 19310
rect 48044 19246 48096 19252
rect 48412 18828 48464 18834
rect 48412 18770 48464 18776
rect 48318 17776 48374 17785
rect 48044 17740 48096 17746
rect 48318 17711 48374 17720
rect 48044 17682 48096 17688
rect 48056 17202 48084 17682
rect 48332 17678 48360 17711
rect 48320 17672 48372 17678
rect 48320 17614 48372 17620
rect 48044 17196 48096 17202
rect 48044 17138 48096 17144
rect 48136 17060 48188 17066
rect 48136 17002 48188 17008
rect 48148 16454 48176 17002
rect 48424 16794 48452 18770
rect 48700 18766 48728 20198
rect 48780 19780 48832 19786
rect 48780 19722 48832 19728
rect 48688 18760 48740 18766
rect 48688 18702 48740 18708
rect 48792 18426 48820 19722
rect 48884 19378 48912 20742
rect 49344 19786 49372 21082
rect 49528 20874 49556 21626
rect 49516 20868 49568 20874
rect 49516 20810 49568 20816
rect 49988 20602 50016 21830
rect 50172 20942 50200 21966
rect 50632 21146 50660 22034
rect 50712 22024 50764 22030
rect 50712 21966 50764 21972
rect 50724 21554 50752 21966
rect 51920 21962 51948 22578
rect 52276 22500 52328 22506
rect 52276 22442 52328 22448
rect 52000 22432 52052 22438
rect 52000 22374 52052 22380
rect 51908 21956 51960 21962
rect 51908 21898 51960 21904
rect 50712 21548 50764 21554
rect 50712 21490 50764 21496
rect 52012 21486 52040 22374
rect 52288 22094 52316 22442
rect 52288 22066 52408 22094
rect 52380 21894 52408 22066
rect 52368 21888 52420 21894
rect 52368 21830 52420 21836
rect 52000 21480 52052 21486
rect 52000 21422 52052 21428
rect 51518 21244 51826 21253
rect 51518 21242 51524 21244
rect 51580 21242 51604 21244
rect 51660 21242 51684 21244
rect 51740 21242 51764 21244
rect 51820 21242 51826 21244
rect 51580 21190 51582 21242
rect 51762 21190 51764 21242
rect 51518 21188 51524 21190
rect 51580 21188 51604 21190
rect 51660 21188 51684 21190
rect 51740 21188 51764 21190
rect 51820 21188 51826 21190
rect 51518 21179 51826 21188
rect 50620 21140 50672 21146
rect 50620 21082 50672 21088
rect 50344 21072 50396 21078
rect 50344 21014 50396 21020
rect 50160 20936 50212 20942
rect 50160 20878 50212 20884
rect 50068 20868 50120 20874
rect 50068 20810 50120 20816
rect 49976 20596 50028 20602
rect 49976 20538 50028 20544
rect 49608 20528 49660 20534
rect 49608 20470 49660 20476
rect 49332 19780 49384 19786
rect 49332 19722 49384 19728
rect 48964 19712 49016 19718
rect 48964 19654 49016 19660
rect 48872 19372 48924 19378
rect 48872 19314 48924 19320
rect 48976 19310 49004 19654
rect 48964 19304 49016 19310
rect 48964 19246 49016 19252
rect 49516 19304 49568 19310
rect 49516 19246 49568 19252
rect 48780 18420 48832 18426
rect 48780 18362 48832 18368
rect 48596 18148 48648 18154
rect 48596 18090 48648 18096
rect 48608 17338 48636 18090
rect 49056 18080 49108 18086
rect 49056 18022 49108 18028
rect 49068 17678 49096 18022
rect 49056 17672 49108 17678
rect 49056 17614 49108 17620
rect 48596 17332 48648 17338
rect 48596 17274 48648 17280
rect 49068 17270 49096 17614
rect 49528 17542 49556 19246
rect 49620 18426 49648 20470
rect 49700 20392 49752 20398
rect 49700 20334 49752 20340
rect 49712 18970 49740 20334
rect 50080 19786 50108 20810
rect 50172 20058 50200 20878
rect 50356 20602 50384 21014
rect 52012 21010 52040 21422
rect 52380 21010 52408 21830
rect 52000 21004 52052 21010
rect 52000 20946 52052 20952
rect 52368 21004 52420 21010
rect 52368 20946 52420 20952
rect 50436 20936 50488 20942
rect 50436 20878 50488 20884
rect 51264 20936 51316 20942
rect 51264 20878 51316 20884
rect 50344 20596 50396 20602
rect 50344 20538 50396 20544
rect 50356 20058 50384 20538
rect 50448 20262 50476 20878
rect 50528 20392 50580 20398
rect 50528 20334 50580 20340
rect 50436 20256 50488 20262
rect 50436 20198 50488 20204
rect 50160 20052 50212 20058
rect 50160 19994 50212 20000
rect 50344 20052 50396 20058
rect 50344 19994 50396 20000
rect 50436 20052 50488 20058
rect 50436 19994 50488 20000
rect 50172 19922 50200 19994
rect 50160 19916 50212 19922
rect 50160 19858 50212 19864
rect 50448 19854 50476 19994
rect 50344 19848 50396 19854
rect 50344 19790 50396 19796
rect 50436 19848 50488 19854
rect 50436 19790 50488 19796
rect 50068 19780 50120 19786
rect 50068 19722 50120 19728
rect 50356 19446 50384 19790
rect 50344 19440 50396 19446
rect 50344 19382 50396 19388
rect 50540 18970 50568 20334
rect 51276 19854 51304 20878
rect 52000 20868 52052 20874
rect 52000 20810 52052 20816
rect 52012 20602 52040 20810
rect 52000 20596 52052 20602
rect 52000 20538 52052 20544
rect 52460 20460 52512 20466
rect 52460 20402 52512 20408
rect 51356 20392 51408 20398
rect 51356 20334 51408 20340
rect 51264 19848 51316 19854
rect 51264 19790 51316 19796
rect 50804 19780 50856 19786
rect 50804 19722 50856 19728
rect 50816 19446 50844 19722
rect 51368 19514 51396 20334
rect 52092 20324 52144 20330
rect 52092 20266 52144 20272
rect 51518 20156 51826 20165
rect 51518 20154 51524 20156
rect 51580 20154 51604 20156
rect 51660 20154 51684 20156
rect 51740 20154 51764 20156
rect 51820 20154 51826 20156
rect 51580 20102 51582 20154
rect 51762 20102 51764 20154
rect 51518 20100 51524 20102
rect 51580 20100 51604 20102
rect 51660 20100 51684 20102
rect 51740 20100 51764 20102
rect 51820 20100 51826 20102
rect 51518 20091 51826 20100
rect 52104 19990 52132 20266
rect 52092 19984 52144 19990
rect 52092 19926 52144 19932
rect 52104 19854 52132 19926
rect 52092 19848 52144 19854
rect 52092 19790 52144 19796
rect 51816 19712 51868 19718
rect 51816 19654 51868 19660
rect 51356 19508 51408 19514
rect 51356 19450 51408 19456
rect 50804 19440 50856 19446
rect 50804 19382 50856 19388
rect 51828 19378 51856 19654
rect 52104 19530 52132 19790
rect 52472 19718 52500 20402
rect 52552 19984 52604 19990
rect 52552 19926 52604 19932
rect 52460 19712 52512 19718
rect 52460 19654 52512 19660
rect 52104 19502 52224 19530
rect 51080 19372 51132 19378
rect 51080 19314 51132 19320
rect 51816 19372 51868 19378
rect 51816 19314 51868 19320
rect 49700 18964 49752 18970
rect 49700 18906 49752 18912
rect 49792 18964 49844 18970
rect 49792 18906 49844 18912
rect 50528 18964 50580 18970
rect 50528 18906 50580 18912
rect 49608 18420 49660 18426
rect 49608 18362 49660 18368
rect 49516 17536 49568 17542
rect 49516 17478 49568 17484
rect 49804 17270 49832 18906
rect 50068 18760 50120 18766
rect 50068 18702 50120 18708
rect 50080 18222 50108 18702
rect 50804 18692 50856 18698
rect 50804 18634 50856 18640
rect 50252 18352 50304 18358
rect 50252 18294 50304 18300
rect 50068 18216 50120 18222
rect 50068 18158 50120 18164
rect 49056 17264 49108 17270
rect 49056 17206 49108 17212
rect 49792 17264 49844 17270
rect 49792 17206 49844 17212
rect 48412 16788 48464 16794
rect 48412 16730 48464 16736
rect 49148 16652 49200 16658
rect 49148 16594 49200 16600
rect 48320 16584 48372 16590
rect 48320 16526 48372 16532
rect 49056 16584 49108 16590
rect 49056 16526 49108 16532
rect 48136 16448 48188 16454
rect 48136 16390 48188 16396
rect 48228 16448 48280 16454
rect 48228 16390 48280 16396
rect 48148 16250 48176 16390
rect 48136 16244 48188 16250
rect 48136 16186 48188 16192
rect 48136 16108 48188 16114
rect 48136 16050 48188 16056
rect 48044 16040 48096 16046
rect 48044 15982 48096 15988
rect 48056 14822 48084 15982
rect 48148 15638 48176 16050
rect 48240 15978 48268 16390
rect 48332 16114 48360 16526
rect 48964 16176 49016 16182
rect 48964 16118 49016 16124
rect 48320 16108 48372 16114
rect 48320 16050 48372 16056
rect 48228 15972 48280 15978
rect 48228 15914 48280 15920
rect 48320 15904 48372 15910
rect 48320 15846 48372 15852
rect 48136 15632 48188 15638
rect 48332 15586 48360 15846
rect 48136 15574 48188 15580
rect 48148 15366 48176 15574
rect 48240 15570 48360 15586
rect 48228 15564 48360 15570
rect 48280 15558 48360 15564
rect 48228 15506 48280 15512
rect 48136 15360 48188 15366
rect 48136 15302 48188 15308
rect 48688 15360 48740 15366
rect 48688 15302 48740 15308
rect 48700 15094 48728 15302
rect 48688 15088 48740 15094
rect 48688 15030 48740 15036
rect 48228 14952 48280 14958
rect 48228 14894 48280 14900
rect 48044 14816 48096 14822
rect 48044 14758 48096 14764
rect 48056 14074 48084 14758
rect 48240 14074 48268 14894
rect 48872 14884 48924 14890
rect 48872 14826 48924 14832
rect 48884 14618 48912 14826
rect 48780 14612 48832 14618
rect 48780 14554 48832 14560
rect 48872 14612 48924 14618
rect 48872 14554 48924 14560
rect 48320 14408 48372 14414
rect 48320 14350 48372 14356
rect 48044 14068 48096 14074
rect 48044 14010 48096 14016
rect 48228 14068 48280 14074
rect 48228 14010 48280 14016
rect 48136 14000 48188 14006
rect 48136 13942 48188 13948
rect 48148 12782 48176 13942
rect 48228 13320 48280 13326
rect 48228 13262 48280 13268
rect 48240 12850 48268 13262
rect 48332 13190 48360 14350
rect 48792 13258 48820 14554
rect 48976 14550 49004 16118
rect 48964 14544 49016 14550
rect 48964 14486 49016 14492
rect 48964 14408 49016 14414
rect 49068 14396 49096 16526
rect 49160 14414 49188 16594
rect 49240 16448 49292 16454
rect 49240 16390 49292 16396
rect 49252 15570 49280 16390
rect 49332 16108 49384 16114
rect 49332 16050 49384 16056
rect 49240 15564 49292 15570
rect 49240 15506 49292 15512
rect 49252 15366 49280 15506
rect 49344 15434 49372 16050
rect 49700 15904 49752 15910
rect 49700 15846 49752 15852
rect 49712 15706 49740 15846
rect 49700 15700 49752 15706
rect 49700 15642 49752 15648
rect 49804 15502 49832 17206
rect 50080 16250 50108 18158
rect 50264 17270 50292 18294
rect 50816 18290 50844 18634
rect 51092 18290 51120 19314
rect 51172 19304 51224 19310
rect 51172 19246 51224 19252
rect 51184 19174 51212 19246
rect 51172 19168 51224 19174
rect 51172 19110 51224 19116
rect 51184 18630 51212 19110
rect 51518 19068 51826 19077
rect 51518 19066 51524 19068
rect 51580 19066 51604 19068
rect 51660 19066 51684 19068
rect 51740 19066 51764 19068
rect 51820 19066 51826 19068
rect 51580 19014 51582 19066
rect 51762 19014 51764 19066
rect 51518 19012 51524 19014
rect 51580 19012 51604 19014
rect 51660 19012 51684 19014
rect 51740 19012 51764 19014
rect 51820 19012 51826 19014
rect 51518 19003 51826 19012
rect 52196 18766 52224 19502
rect 52472 18834 52500 19654
rect 52564 19242 52592 19926
rect 52552 19236 52604 19242
rect 52552 19178 52604 19184
rect 52460 18828 52512 18834
rect 52460 18770 52512 18776
rect 52184 18760 52236 18766
rect 52184 18702 52236 18708
rect 52368 18692 52420 18698
rect 52564 18680 52592 19178
rect 52656 18902 52684 32710
rect 56612 31142 56640 33390
rect 57520 33312 57572 33318
rect 57520 33254 57572 33260
rect 56600 31136 56652 31142
rect 56600 31078 56652 31084
rect 56600 23724 56652 23730
rect 56600 23666 56652 23672
rect 55128 22024 55180 22030
rect 56612 22001 56640 23666
rect 55128 21966 55180 21972
rect 56598 21992 56654 22001
rect 53104 21548 53156 21554
rect 53104 21490 53156 21496
rect 52828 21344 52880 21350
rect 52828 21286 52880 21292
rect 52840 20602 52868 21286
rect 52828 20596 52880 20602
rect 52828 20538 52880 20544
rect 52840 19922 52868 20538
rect 52920 20256 52972 20262
rect 52920 20198 52972 20204
rect 52828 19916 52880 19922
rect 52828 19858 52880 19864
rect 52932 19394 52960 20198
rect 53012 19916 53064 19922
rect 53012 19858 53064 19864
rect 53024 19514 53052 19858
rect 53116 19854 53144 21490
rect 55140 21486 55168 21966
rect 56598 21927 56654 21936
rect 55588 21888 55640 21894
rect 55588 21830 55640 21836
rect 54300 21480 54352 21486
rect 54300 21422 54352 21428
rect 55128 21480 55180 21486
rect 55128 21422 55180 21428
rect 53656 21004 53708 21010
rect 53656 20946 53708 20952
rect 53288 20936 53340 20942
rect 53288 20878 53340 20884
rect 53300 20806 53328 20878
rect 53288 20800 53340 20806
rect 53288 20742 53340 20748
rect 53472 20800 53524 20806
rect 53472 20742 53524 20748
rect 53300 20602 53328 20742
rect 53288 20596 53340 20602
rect 53288 20538 53340 20544
rect 53484 20534 53512 20742
rect 53472 20528 53524 20534
rect 53472 20470 53524 20476
rect 53196 20052 53248 20058
rect 53196 19994 53248 20000
rect 53104 19848 53156 19854
rect 53104 19790 53156 19796
rect 53012 19508 53064 19514
rect 53012 19450 53064 19456
rect 52932 19378 53052 19394
rect 52828 19372 52880 19378
rect 52932 19372 53064 19378
rect 52932 19366 53012 19372
rect 52828 19314 52880 19320
rect 53012 19314 53064 19320
rect 52840 18970 52868 19314
rect 53208 18970 53236 19994
rect 53668 19990 53696 20946
rect 54116 20936 54168 20942
rect 54116 20878 54168 20884
rect 54128 20602 54156 20878
rect 54116 20596 54168 20602
rect 54116 20538 54168 20544
rect 53748 20392 53800 20398
rect 53748 20334 53800 20340
rect 53656 19984 53708 19990
rect 53656 19926 53708 19932
rect 53760 19854 53788 20334
rect 53840 20324 53892 20330
rect 53840 20266 53892 20272
rect 53656 19848 53708 19854
rect 53656 19790 53708 19796
rect 53748 19848 53800 19854
rect 53748 19790 53800 19796
rect 53288 19712 53340 19718
rect 53288 19654 53340 19660
rect 53300 19242 53328 19654
rect 53668 19514 53696 19790
rect 53852 19786 53880 20266
rect 53840 19780 53892 19786
rect 53840 19722 53892 19728
rect 53656 19508 53708 19514
rect 53656 19450 53708 19456
rect 53288 19236 53340 19242
rect 53288 19178 53340 19184
rect 53852 19174 53880 19722
rect 54312 19378 54340 21422
rect 55496 21344 55548 21350
rect 55496 21286 55548 21292
rect 55508 21146 55536 21286
rect 55496 21140 55548 21146
rect 55496 21082 55548 21088
rect 55508 20942 55536 21082
rect 55496 20936 55548 20942
rect 55496 20878 55548 20884
rect 55220 20256 55272 20262
rect 55220 20198 55272 20204
rect 54760 19848 54812 19854
rect 54760 19790 54812 19796
rect 53932 19372 53984 19378
rect 53932 19314 53984 19320
rect 54300 19372 54352 19378
rect 54300 19314 54352 19320
rect 53840 19168 53892 19174
rect 53840 19110 53892 19116
rect 52828 18964 52880 18970
rect 52828 18906 52880 18912
rect 53196 18964 53248 18970
rect 53196 18906 53248 18912
rect 52644 18896 52696 18902
rect 52644 18838 52696 18844
rect 52920 18828 52972 18834
rect 52920 18770 52972 18776
rect 53196 18828 53248 18834
rect 53196 18770 53248 18776
rect 52564 18652 52684 18680
rect 52368 18634 52420 18640
rect 51172 18624 51224 18630
rect 51172 18566 51224 18572
rect 50804 18284 50856 18290
rect 50804 18226 50856 18232
rect 51080 18284 51132 18290
rect 51080 18226 51132 18232
rect 52000 18284 52052 18290
rect 52000 18226 52052 18232
rect 52184 18284 52236 18290
rect 52184 18226 52236 18232
rect 50528 18216 50580 18222
rect 50528 18158 50580 18164
rect 50436 18080 50488 18086
rect 50436 18022 50488 18028
rect 50448 17746 50476 18022
rect 50540 17882 50568 18158
rect 50528 17876 50580 17882
rect 50528 17818 50580 17824
rect 50436 17740 50488 17746
rect 50436 17682 50488 17688
rect 50252 17264 50304 17270
rect 50252 17206 50304 17212
rect 50160 17128 50212 17134
rect 50160 17070 50212 17076
rect 50172 16794 50200 17070
rect 50160 16788 50212 16794
rect 50160 16730 50212 16736
rect 50068 16244 50120 16250
rect 50068 16186 50120 16192
rect 49792 15496 49844 15502
rect 49792 15438 49844 15444
rect 49332 15428 49384 15434
rect 49332 15370 49384 15376
rect 49240 15360 49292 15366
rect 49240 15302 49292 15308
rect 49804 14958 49832 15438
rect 49976 15360 50028 15366
rect 49976 15302 50028 15308
rect 49792 14952 49844 14958
rect 49792 14894 49844 14900
rect 49700 14816 49752 14822
rect 49700 14758 49752 14764
rect 49016 14368 49096 14396
rect 49148 14408 49200 14414
rect 48964 14350 49016 14356
rect 49200 14368 49280 14396
rect 49148 14350 49200 14356
rect 48976 14278 49004 14350
rect 48964 14272 49016 14278
rect 48964 14214 49016 14220
rect 49252 14074 49280 14368
rect 49240 14068 49292 14074
rect 49240 14010 49292 14016
rect 49148 13728 49200 13734
rect 49148 13670 49200 13676
rect 48780 13252 48832 13258
rect 48780 13194 48832 13200
rect 48320 13184 48372 13190
rect 48320 13126 48372 13132
rect 48792 12986 48820 13194
rect 48780 12980 48832 12986
rect 48780 12922 48832 12928
rect 48228 12844 48280 12850
rect 48228 12786 48280 12792
rect 48136 12776 48188 12782
rect 48136 12718 48188 12724
rect 48148 12186 48176 12718
rect 48240 12442 48268 12786
rect 49160 12782 49188 13670
rect 49332 13184 49384 13190
rect 49332 13126 49384 13132
rect 49344 12850 49372 13126
rect 49332 12844 49384 12850
rect 49332 12786 49384 12792
rect 49148 12776 49200 12782
rect 49148 12718 49200 12724
rect 48688 12708 48740 12714
rect 48688 12650 48740 12656
rect 48412 12640 48464 12646
rect 48412 12582 48464 12588
rect 48228 12436 48280 12442
rect 48228 12378 48280 12384
rect 48148 12170 48268 12186
rect 48148 12164 48280 12170
rect 48148 12158 48228 12164
rect 48228 12106 48280 12112
rect 48240 11830 48268 12106
rect 48320 11892 48372 11898
rect 48320 11834 48372 11840
rect 48228 11824 48280 11830
rect 48228 11766 48280 11772
rect 48136 11756 48188 11762
rect 47964 11716 48136 11744
rect 48136 11698 48188 11704
rect 47860 11552 47912 11558
rect 47860 11494 47912 11500
rect 47872 11150 47900 11494
rect 47860 11144 47912 11150
rect 47860 11086 47912 11092
rect 48044 11144 48096 11150
rect 48044 11086 48096 11092
rect 48056 10742 48084 11086
rect 48148 11014 48176 11698
rect 48228 11212 48280 11218
rect 48332 11200 48360 11834
rect 48280 11172 48360 11200
rect 48228 11154 48280 11160
rect 48136 11008 48188 11014
rect 48136 10950 48188 10956
rect 48044 10736 48096 10742
rect 48044 10678 48096 10684
rect 48056 10470 48084 10678
rect 48148 10606 48176 10950
rect 48136 10600 48188 10606
rect 48136 10542 48188 10548
rect 48044 10464 48096 10470
rect 48044 10406 48096 10412
rect 48056 10266 48084 10406
rect 48044 10260 48096 10266
rect 48044 10202 48096 10208
rect 48228 9580 48280 9586
rect 48228 9522 48280 9528
rect 48240 9178 48268 9522
rect 48332 9518 48360 11172
rect 48320 9512 48372 9518
rect 48320 9454 48372 9460
rect 48228 9172 48280 9178
rect 48228 9114 48280 9120
rect 46388 8832 46440 8838
rect 46388 8774 46440 8780
rect 47676 8832 47728 8838
rect 47676 8774 47728 8780
rect 46204 8628 46256 8634
rect 46204 8570 46256 8576
rect 46400 8498 46428 8774
rect 46388 8492 46440 8498
rect 46388 8434 46440 8440
rect 46572 8492 46624 8498
rect 46572 8434 46624 8440
rect 47308 8492 47360 8498
rect 47308 8434 47360 8440
rect 46400 8265 46428 8434
rect 46386 8256 46442 8265
rect 46386 8191 46442 8200
rect 46400 7954 46428 8191
rect 46388 7948 46440 7954
rect 46440 7908 46520 7936
rect 46388 7890 46440 7896
rect 46296 7880 46348 7886
rect 46296 7822 46348 7828
rect 46308 7546 46336 7822
rect 46388 7744 46440 7750
rect 46388 7686 46440 7692
rect 46296 7540 46348 7546
rect 46296 7482 46348 7488
rect 45928 7404 45980 7410
rect 45928 7346 45980 7352
rect 45940 6798 45968 7346
rect 46400 7002 46428 7686
rect 46492 7002 46520 7908
rect 46584 7546 46612 8434
rect 47320 8090 47348 8434
rect 47308 8084 47360 8090
rect 47308 8026 47360 8032
rect 47124 7812 47176 7818
rect 47124 7754 47176 7760
rect 46572 7540 46624 7546
rect 46572 7482 46624 7488
rect 47136 7478 47164 7754
rect 47124 7472 47176 7478
rect 47124 7414 47176 7420
rect 46388 6996 46440 7002
rect 46388 6938 46440 6944
rect 46480 6996 46532 7002
rect 46480 6938 46532 6944
rect 45560 6792 45612 6798
rect 45560 6734 45612 6740
rect 45928 6792 45980 6798
rect 45928 6734 45980 6740
rect 44732 6724 44784 6730
rect 44732 6666 44784 6672
rect 44294 6556 44602 6565
rect 44294 6554 44300 6556
rect 44356 6554 44380 6556
rect 44436 6554 44460 6556
rect 44516 6554 44540 6556
rect 44596 6554 44602 6556
rect 44356 6502 44358 6554
rect 44538 6502 44540 6554
rect 44294 6500 44300 6502
rect 44356 6500 44380 6502
rect 44436 6500 44460 6502
rect 44516 6500 44540 6502
rect 44596 6500 44602 6502
rect 44294 6491 44602 6500
rect 45940 6458 45968 6734
rect 45928 6452 45980 6458
rect 45928 6394 45980 6400
rect 44294 5468 44602 5477
rect 44294 5466 44300 5468
rect 44356 5466 44380 5468
rect 44436 5466 44460 5468
rect 44516 5466 44540 5468
rect 44596 5466 44602 5468
rect 44356 5414 44358 5466
rect 44538 5414 44540 5466
rect 44294 5412 44300 5414
rect 44356 5412 44380 5414
rect 44436 5412 44460 5414
rect 44516 5412 44540 5414
rect 44596 5412 44602 5414
rect 44294 5403 44602 5412
rect 44294 4380 44602 4389
rect 44294 4378 44300 4380
rect 44356 4378 44380 4380
rect 44436 4378 44460 4380
rect 44516 4378 44540 4380
rect 44596 4378 44602 4380
rect 44356 4326 44358 4378
rect 44538 4326 44540 4378
rect 44294 4324 44300 4326
rect 44356 4324 44380 4326
rect 44436 4324 44460 4326
rect 44516 4324 44540 4326
rect 44596 4324 44602 4326
rect 44294 4315 44602 4324
rect 44294 3292 44602 3301
rect 44294 3290 44300 3292
rect 44356 3290 44380 3292
rect 44436 3290 44460 3292
rect 44516 3290 44540 3292
rect 44596 3290 44602 3292
rect 44356 3238 44358 3290
rect 44538 3238 44540 3290
rect 44294 3236 44300 3238
rect 44356 3236 44380 3238
rect 44436 3236 44460 3238
rect 44516 3236 44540 3238
rect 44596 3236 44602 3238
rect 44294 3227 44602 3236
rect 44180 3188 44232 3194
rect 44180 3130 44232 3136
rect 48424 2446 48452 12582
rect 48700 12306 48728 12650
rect 49712 12306 49740 14758
rect 49988 13870 50016 15302
rect 50264 15094 50292 17206
rect 50620 16652 50672 16658
rect 50620 16594 50672 16600
rect 50632 15473 50660 16594
rect 51092 15502 51120 18226
rect 51518 17980 51826 17989
rect 51518 17978 51524 17980
rect 51580 17978 51604 17980
rect 51660 17978 51684 17980
rect 51740 17978 51764 17980
rect 51820 17978 51826 17980
rect 51580 17926 51582 17978
rect 51762 17926 51764 17978
rect 51518 17924 51524 17926
rect 51580 17924 51604 17926
rect 51660 17924 51684 17926
rect 51740 17924 51764 17926
rect 51820 17924 51826 17926
rect 51518 17915 51826 17924
rect 51906 17912 51962 17921
rect 51906 17847 51962 17856
rect 51816 17672 51868 17678
rect 51816 17614 51868 17620
rect 51828 17338 51856 17614
rect 51816 17332 51868 17338
rect 51816 17274 51868 17280
rect 51920 17202 51948 17847
rect 51908 17196 51960 17202
rect 51908 17138 51960 17144
rect 51448 17060 51500 17066
rect 51448 17002 51500 17008
rect 51356 16992 51408 16998
rect 51356 16934 51408 16940
rect 51368 16726 51396 16934
rect 51356 16720 51408 16726
rect 51356 16662 51408 16668
rect 51368 16114 51396 16662
rect 51460 16658 51488 17002
rect 51518 16892 51826 16901
rect 51518 16890 51524 16892
rect 51580 16890 51604 16892
rect 51660 16890 51684 16892
rect 51740 16890 51764 16892
rect 51820 16890 51826 16892
rect 51580 16838 51582 16890
rect 51762 16838 51764 16890
rect 51518 16836 51524 16838
rect 51580 16836 51604 16838
rect 51660 16836 51684 16838
rect 51740 16836 51764 16838
rect 51820 16836 51826 16838
rect 51518 16827 51826 16836
rect 51448 16652 51500 16658
rect 51448 16594 51500 16600
rect 52012 16590 52040 18226
rect 52196 17882 52224 18226
rect 52184 17876 52236 17882
rect 52184 17818 52236 17824
rect 52380 17746 52408 18634
rect 52368 17740 52420 17746
rect 52368 17682 52420 17688
rect 52460 17672 52512 17678
rect 52460 17614 52512 17620
rect 52184 17604 52236 17610
rect 52184 17546 52236 17552
rect 52196 17066 52224 17546
rect 52368 17128 52420 17134
rect 52368 17070 52420 17076
rect 52184 17060 52236 17066
rect 52184 17002 52236 17008
rect 52000 16584 52052 16590
rect 52000 16526 52052 16532
rect 52380 16504 52408 17070
rect 52472 16794 52500 17614
rect 52552 17196 52604 17202
rect 52552 17138 52604 17144
rect 52564 16998 52592 17138
rect 52552 16992 52604 16998
rect 52552 16934 52604 16940
rect 52460 16788 52512 16794
rect 52460 16730 52512 16736
rect 52460 16516 52512 16522
rect 52380 16476 52460 16504
rect 52460 16458 52512 16464
rect 52472 16250 52500 16458
rect 52656 16402 52684 18652
rect 52736 18352 52788 18358
rect 52736 18294 52788 18300
rect 52748 17610 52776 18294
rect 52828 18284 52880 18290
rect 52828 18226 52880 18232
rect 52736 17604 52788 17610
rect 52736 17546 52788 17552
rect 52748 17202 52776 17546
rect 52736 17196 52788 17202
rect 52736 17138 52788 17144
rect 52736 16992 52788 16998
rect 52736 16934 52788 16940
rect 52748 16538 52776 16934
rect 52840 16726 52868 18226
rect 52932 17678 52960 18770
rect 53208 18222 53236 18770
rect 53288 18284 53340 18290
rect 53288 18226 53340 18232
rect 53196 18216 53248 18222
rect 53196 18158 53248 18164
rect 53012 18148 53064 18154
rect 53012 18090 53064 18096
rect 52920 17672 52972 17678
rect 52920 17614 52972 17620
rect 53024 17542 53052 18090
rect 53208 17882 53236 18158
rect 53196 17876 53248 17882
rect 53196 17818 53248 17824
rect 53300 17542 53328 18226
rect 53472 18148 53524 18154
rect 53472 18090 53524 18096
rect 53484 17610 53512 18090
rect 53564 18080 53616 18086
rect 53564 18022 53616 18028
rect 53840 18080 53892 18086
rect 53840 18022 53892 18028
rect 53472 17604 53524 17610
rect 53472 17546 53524 17552
rect 53012 17536 53064 17542
rect 53012 17478 53064 17484
rect 53288 17536 53340 17542
rect 53288 17478 53340 17484
rect 52920 17264 52972 17270
rect 52920 17206 52972 17212
rect 52828 16720 52880 16726
rect 52828 16662 52880 16668
rect 52748 16510 52868 16538
rect 52840 16454 52868 16510
rect 52564 16374 52684 16402
rect 52736 16448 52788 16454
rect 52736 16390 52788 16396
rect 52828 16448 52880 16454
rect 52828 16390 52880 16396
rect 52460 16244 52512 16250
rect 52460 16186 52512 16192
rect 51356 16108 51408 16114
rect 51356 16050 51408 16056
rect 52564 16046 52592 16374
rect 52748 16114 52776 16390
rect 52736 16108 52788 16114
rect 52736 16050 52788 16056
rect 52552 16040 52604 16046
rect 51170 16008 51226 16017
rect 52552 15982 52604 15988
rect 51170 15943 51226 15952
rect 51184 15706 51212 15943
rect 51264 15904 51316 15910
rect 51264 15846 51316 15852
rect 51172 15700 51224 15706
rect 51172 15642 51224 15648
rect 51276 15502 51304 15846
rect 51518 15804 51826 15813
rect 51518 15802 51524 15804
rect 51580 15802 51604 15804
rect 51660 15802 51684 15804
rect 51740 15802 51764 15804
rect 51820 15802 51826 15804
rect 51580 15750 51582 15802
rect 51762 15750 51764 15802
rect 51518 15748 51524 15750
rect 51580 15748 51604 15750
rect 51660 15748 51684 15750
rect 51740 15748 51764 15750
rect 51820 15748 51826 15750
rect 51518 15739 51826 15748
rect 51080 15496 51132 15502
rect 50618 15464 50674 15473
rect 50986 15464 51042 15473
rect 50618 15399 50674 15408
rect 50712 15428 50764 15434
rect 51080 15438 51132 15444
rect 51264 15496 51316 15502
rect 51264 15438 51316 15444
rect 52184 15496 52236 15502
rect 52184 15438 52236 15444
rect 50986 15399 51042 15408
rect 50712 15370 50764 15376
rect 50724 15162 50752 15370
rect 50712 15156 50764 15162
rect 50712 15098 50764 15104
rect 50252 15088 50304 15094
rect 50252 15030 50304 15036
rect 50896 14476 50948 14482
rect 50896 14418 50948 14424
rect 50908 14278 50936 14418
rect 50344 14272 50396 14278
rect 50344 14214 50396 14220
rect 50712 14272 50764 14278
rect 50712 14214 50764 14220
rect 50896 14272 50948 14278
rect 50896 14214 50948 14220
rect 49976 13864 50028 13870
rect 49976 13806 50028 13812
rect 49792 13252 49844 13258
rect 49792 13194 49844 13200
rect 48688 12300 48740 12306
rect 48688 12242 48740 12248
rect 49700 12300 49752 12306
rect 49700 12242 49752 12248
rect 49516 11892 49568 11898
rect 49516 11834 49568 11840
rect 48504 11688 48556 11694
rect 48504 11630 48556 11636
rect 48516 11286 48544 11630
rect 48964 11552 49016 11558
rect 48964 11494 49016 11500
rect 48504 11280 48556 11286
rect 48504 11222 48556 11228
rect 48976 10674 49004 11494
rect 49528 10674 49556 11834
rect 49700 11756 49752 11762
rect 49700 11698 49752 11704
rect 49712 11150 49740 11698
rect 49804 11150 49832 13194
rect 49988 12442 50016 13806
rect 50356 13326 50384 14214
rect 50620 14068 50672 14074
rect 50620 14010 50672 14016
rect 50632 13462 50660 14010
rect 50620 13456 50672 13462
rect 50620 13398 50672 13404
rect 50344 13320 50396 13326
rect 50344 13262 50396 13268
rect 50252 12912 50304 12918
rect 50252 12854 50304 12860
rect 49976 12436 50028 12442
rect 49976 12378 50028 12384
rect 50264 11558 50292 12854
rect 50356 12850 50384 13262
rect 50436 12980 50488 12986
rect 50724 12968 50752 14214
rect 50908 14006 50936 14214
rect 50896 14000 50948 14006
rect 50896 13942 50948 13948
rect 50804 13320 50856 13326
rect 50804 13262 50856 13268
rect 50488 12940 50752 12968
rect 50436 12922 50488 12928
rect 50344 12844 50396 12850
rect 50344 12786 50396 12792
rect 50436 12232 50488 12238
rect 50724 12220 50752 12940
rect 50816 12782 50844 13262
rect 50804 12776 50856 12782
rect 50804 12718 50856 12724
rect 50816 12442 50844 12718
rect 50804 12436 50856 12442
rect 50804 12378 50856 12384
rect 50804 12232 50856 12238
rect 50724 12192 50804 12220
rect 50436 12174 50488 12180
rect 50804 12174 50856 12180
rect 50448 11694 50476 12174
rect 50896 11756 50948 11762
rect 50896 11698 50948 11704
rect 50436 11688 50488 11694
rect 50436 11630 50488 11636
rect 50252 11552 50304 11558
rect 50252 11494 50304 11500
rect 49700 11144 49752 11150
rect 49700 11086 49752 11092
rect 49792 11144 49844 11150
rect 49792 11086 49844 11092
rect 49712 10742 49740 11086
rect 49700 10736 49752 10742
rect 49700 10678 49752 10684
rect 48964 10668 49016 10674
rect 48964 10610 49016 10616
rect 49516 10668 49568 10674
rect 49516 10610 49568 10616
rect 49804 9722 49832 11086
rect 49792 9716 49844 9722
rect 49792 9658 49844 9664
rect 50264 9586 50292 11494
rect 50908 11082 50936 11698
rect 50896 11076 50948 11082
rect 50896 11018 50948 11024
rect 50252 9580 50304 9586
rect 50252 9522 50304 9528
rect 51000 9178 51028 15399
rect 51092 12434 51120 15438
rect 51908 15360 51960 15366
rect 51908 15302 51960 15308
rect 51356 15020 51408 15026
rect 51356 14962 51408 14968
rect 51264 14816 51316 14822
rect 51264 14758 51316 14764
rect 51172 14340 51224 14346
rect 51172 14282 51224 14288
rect 51184 13938 51212 14282
rect 51276 14074 51304 14758
rect 51368 14414 51396 14962
rect 51448 14952 51500 14958
rect 51448 14894 51500 14900
rect 51460 14414 51488 14894
rect 51518 14716 51826 14725
rect 51518 14714 51524 14716
rect 51580 14714 51604 14716
rect 51660 14714 51684 14716
rect 51740 14714 51764 14716
rect 51820 14714 51826 14716
rect 51580 14662 51582 14714
rect 51762 14662 51764 14714
rect 51518 14660 51524 14662
rect 51580 14660 51604 14662
rect 51660 14660 51684 14662
rect 51740 14660 51764 14662
rect 51820 14660 51826 14662
rect 51518 14651 51826 14660
rect 51920 14482 51948 15302
rect 52196 15162 52224 15438
rect 52184 15156 52236 15162
rect 52184 15098 52236 15104
rect 51908 14476 51960 14482
rect 51908 14418 51960 14424
rect 51356 14408 51408 14414
rect 51356 14350 51408 14356
rect 51448 14408 51500 14414
rect 51448 14350 51500 14356
rect 51908 14272 51960 14278
rect 51908 14214 51960 14220
rect 51264 14068 51316 14074
rect 51264 14010 51316 14016
rect 51172 13932 51224 13938
rect 51172 13874 51224 13880
rect 51356 13864 51408 13870
rect 51356 13806 51408 13812
rect 51368 13326 51396 13806
rect 51518 13628 51826 13637
rect 51518 13626 51524 13628
rect 51580 13626 51604 13628
rect 51660 13626 51684 13628
rect 51740 13626 51764 13628
rect 51820 13626 51826 13628
rect 51580 13574 51582 13626
rect 51762 13574 51764 13626
rect 51518 13572 51524 13574
rect 51580 13572 51604 13574
rect 51660 13572 51684 13574
rect 51740 13572 51764 13574
rect 51820 13572 51826 13574
rect 51518 13563 51826 13572
rect 51920 13394 51948 14214
rect 52196 13938 52224 15098
rect 52368 14544 52420 14550
rect 52368 14486 52420 14492
rect 52184 13932 52236 13938
rect 52184 13874 52236 13880
rect 51908 13388 51960 13394
rect 51908 13330 51960 13336
rect 51356 13320 51408 13326
rect 51356 13262 51408 13268
rect 51908 12912 51960 12918
rect 51908 12854 51960 12860
rect 51518 12540 51826 12549
rect 51518 12538 51524 12540
rect 51580 12538 51604 12540
rect 51660 12538 51684 12540
rect 51740 12538 51764 12540
rect 51820 12538 51826 12540
rect 51580 12486 51582 12538
rect 51762 12486 51764 12538
rect 51518 12484 51524 12486
rect 51580 12484 51604 12486
rect 51660 12484 51684 12486
rect 51740 12484 51764 12486
rect 51820 12484 51826 12486
rect 51518 12475 51826 12484
rect 51920 12442 51948 12854
rect 52380 12646 52408 14486
rect 52368 12640 52420 12646
rect 52368 12582 52420 12588
rect 51908 12436 51960 12442
rect 51092 12406 51212 12434
rect 51080 12096 51132 12102
rect 51184 12084 51212 12406
rect 51908 12378 51960 12384
rect 52564 12170 52592 15982
rect 52748 15434 52776 16050
rect 52828 15564 52880 15570
rect 52828 15506 52880 15512
rect 52840 15473 52868 15506
rect 52826 15464 52882 15473
rect 52736 15428 52788 15434
rect 52826 15399 52882 15408
rect 52736 15370 52788 15376
rect 52828 15360 52880 15366
rect 52828 15302 52880 15308
rect 52840 15094 52868 15302
rect 52828 15088 52880 15094
rect 52828 15030 52880 15036
rect 52932 14618 52960 17206
rect 52920 14612 52972 14618
rect 52920 14554 52972 14560
rect 52920 14340 52972 14346
rect 52920 14282 52972 14288
rect 52932 13530 52960 14282
rect 52920 13524 52972 13530
rect 52920 13466 52972 13472
rect 53024 12850 53052 17478
rect 53484 17338 53512 17546
rect 53576 17338 53604 18022
rect 53852 17921 53880 18022
rect 53838 17912 53894 17921
rect 53944 17882 53972 19314
rect 54772 18834 54800 19790
rect 54760 18828 54812 18834
rect 54760 18770 54812 18776
rect 54208 18624 54260 18630
rect 54208 18566 54260 18572
rect 54116 18216 54168 18222
rect 54116 18158 54168 18164
rect 53838 17847 53894 17856
rect 53932 17876 53984 17882
rect 53932 17818 53984 17824
rect 54128 17678 54156 18158
rect 54116 17672 54168 17678
rect 54116 17614 54168 17620
rect 53472 17332 53524 17338
rect 53472 17274 53524 17280
rect 53564 17332 53616 17338
rect 53564 17274 53616 17280
rect 53196 16992 53248 16998
rect 53196 16934 53248 16940
rect 53208 16522 53236 16934
rect 53380 16720 53432 16726
rect 53380 16662 53432 16668
rect 53288 16584 53340 16590
rect 53288 16526 53340 16532
rect 53196 16516 53248 16522
rect 53196 16458 53248 16464
rect 53196 15972 53248 15978
rect 53196 15914 53248 15920
rect 53208 15434 53236 15914
rect 53196 15428 53248 15434
rect 53196 15370 53248 15376
rect 53208 15042 53236 15370
rect 53116 15026 53236 15042
rect 53300 15026 53328 16526
rect 53392 16182 53420 16662
rect 53380 16176 53432 16182
rect 53380 16118 53432 16124
rect 53380 15700 53432 15706
rect 53380 15642 53432 15648
rect 53104 15020 53236 15026
rect 53156 15014 53236 15020
rect 53104 14962 53156 14968
rect 53208 14482 53236 15014
rect 53288 15020 53340 15026
rect 53288 14962 53340 14968
rect 53196 14476 53248 14482
rect 53196 14418 53248 14424
rect 53300 14414 53328 14962
rect 53392 14822 53420 15642
rect 53484 15042 53512 17274
rect 54220 17134 54248 18566
rect 54300 17740 54352 17746
rect 54300 17682 54352 17688
rect 54208 17128 54260 17134
rect 54208 17070 54260 17076
rect 53932 17060 53984 17066
rect 53932 17002 53984 17008
rect 53944 16590 53972 17002
rect 54312 16794 54340 17682
rect 54772 17678 54800 18770
rect 54760 17672 54812 17678
rect 54760 17614 54812 17620
rect 54392 17604 54444 17610
rect 54392 17546 54444 17552
rect 54300 16788 54352 16794
rect 54300 16730 54352 16736
rect 54404 16658 54432 17546
rect 55232 17202 55260 20198
rect 55600 19922 55628 21830
rect 56692 21548 56744 21554
rect 56692 21490 56744 21496
rect 55772 21480 55824 21486
rect 55772 21422 55824 21428
rect 55784 21146 55812 21422
rect 55772 21140 55824 21146
rect 55772 21082 55824 21088
rect 56704 20942 56732 21490
rect 56692 20936 56744 20942
rect 56692 20878 56744 20884
rect 57336 20868 57388 20874
rect 57336 20810 57388 20816
rect 55588 19916 55640 19922
rect 55588 19858 55640 19864
rect 56324 19916 56376 19922
rect 56324 19858 56376 19864
rect 56232 18216 56284 18222
rect 56232 18158 56284 18164
rect 55956 18080 56008 18086
rect 55956 18022 56008 18028
rect 55968 17270 55996 18022
rect 56244 17338 56272 18158
rect 56336 17746 56364 19858
rect 57348 19786 57376 20810
rect 57336 19780 57388 19786
rect 57336 19722 57388 19728
rect 57348 19446 57376 19722
rect 57336 19440 57388 19446
rect 57336 19382 57388 19388
rect 57348 18766 57376 19382
rect 57336 18760 57388 18766
rect 57336 18702 57388 18708
rect 56416 18284 56468 18290
rect 56416 18226 56468 18232
rect 56428 17882 56456 18226
rect 56692 18148 56744 18154
rect 56692 18090 56744 18096
rect 56416 17876 56468 17882
rect 56416 17818 56468 17824
rect 56324 17740 56376 17746
rect 56324 17682 56376 17688
rect 56232 17332 56284 17338
rect 56232 17274 56284 17280
rect 55956 17264 56008 17270
rect 55956 17206 56008 17212
rect 55036 17196 55088 17202
rect 55036 17138 55088 17144
rect 55220 17196 55272 17202
rect 55220 17138 55272 17144
rect 54392 16652 54444 16658
rect 54392 16594 54444 16600
rect 53932 16584 53984 16590
rect 53932 16526 53984 16532
rect 54116 16448 54168 16454
rect 54116 16390 54168 16396
rect 53564 16176 53616 16182
rect 53564 16118 53616 16124
rect 53576 15434 53604 16118
rect 54128 16114 54156 16390
rect 54208 16244 54260 16250
rect 54208 16186 54260 16192
rect 54116 16108 54168 16114
rect 54116 16050 54168 16056
rect 53748 15904 53800 15910
rect 53748 15846 53800 15852
rect 53564 15428 53616 15434
rect 53564 15370 53616 15376
rect 53656 15360 53708 15366
rect 53656 15302 53708 15308
rect 53484 15014 53604 15042
rect 53472 14952 53524 14958
rect 53472 14894 53524 14900
rect 53380 14816 53432 14822
rect 53380 14758 53432 14764
rect 53392 14414 53420 14758
rect 53288 14408 53340 14414
rect 53288 14350 53340 14356
rect 53380 14408 53432 14414
rect 53380 14350 53432 14356
rect 53484 14346 53512 14894
rect 53472 14340 53524 14346
rect 53472 14282 53524 14288
rect 53484 14006 53512 14282
rect 53472 14000 53524 14006
rect 53472 13942 53524 13948
rect 53196 13932 53248 13938
rect 53196 13874 53248 13880
rect 53208 13258 53236 13874
rect 53380 13388 53432 13394
rect 53380 13330 53432 13336
rect 53196 13252 53248 13258
rect 53196 13194 53248 13200
rect 53208 12986 53236 13194
rect 53392 12986 53420 13330
rect 53576 13326 53604 15014
rect 53668 14414 53696 15302
rect 53760 14958 53788 15846
rect 54128 15502 54156 16050
rect 54220 15502 54248 16186
rect 53840 15496 53892 15502
rect 53840 15438 53892 15444
rect 54116 15496 54168 15502
rect 54116 15438 54168 15444
rect 54208 15496 54260 15502
rect 54208 15438 54260 15444
rect 53748 14952 53800 14958
rect 53748 14894 53800 14900
rect 53656 14408 53708 14414
rect 53656 14350 53708 14356
rect 53852 14074 53880 15438
rect 54024 14408 54076 14414
rect 54024 14350 54076 14356
rect 53840 14068 53892 14074
rect 53840 14010 53892 14016
rect 54036 13938 54064 14350
rect 54024 13932 54076 13938
rect 54024 13874 54076 13880
rect 54208 13932 54260 13938
rect 54208 13874 54260 13880
rect 54220 13802 54248 13874
rect 54208 13796 54260 13802
rect 54208 13738 54260 13744
rect 53564 13320 53616 13326
rect 53564 13262 53616 13268
rect 53576 12986 53604 13262
rect 53196 12980 53248 12986
rect 53196 12922 53248 12928
rect 53380 12980 53432 12986
rect 53380 12922 53432 12928
rect 53564 12980 53616 12986
rect 53564 12922 53616 12928
rect 53012 12844 53064 12850
rect 53012 12786 53064 12792
rect 53024 12442 53052 12786
rect 53380 12776 53432 12782
rect 53380 12718 53432 12724
rect 53012 12436 53064 12442
rect 53012 12378 53064 12384
rect 53392 12170 53420 12718
rect 53576 12434 53604 12922
rect 53932 12708 53984 12714
rect 53932 12650 53984 12656
rect 53484 12406 53604 12434
rect 53484 12306 53512 12406
rect 53472 12300 53524 12306
rect 53472 12242 53524 12248
rect 52552 12164 52604 12170
rect 52552 12106 52604 12112
rect 53380 12164 53432 12170
rect 53380 12106 53432 12112
rect 53840 12164 53892 12170
rect 53840 12106 53892 12112
rect 51132 12056 51212 12084
rect 53012 12096 53064 12102
rect 51080 12038 51132 12044
rect 53012 12038 53064 12044
rect 51092 11694 51120 12038
rect 53024 11694 53052 12038
rect 53288 11756 53340 11762
rect 53852 11744 53880 12106
rect 53944 11898 53972 12650
rect 54404 12442 54432 16594
rect 54760 16108 54812 16114
rect 54760 16050 54812 16056
rect 54944 16108 54996 16114
rect 54944 16050 54996 16056
rect 54772 15706 54800 16050
rect 54760 15700 54812 15706
rect 54760 15642 54812 15648
rect 54956 15638 54984 16050
rect 55048 16046 55076 17138
rect 55232 16590 55260 17138
rect 56336 16658 56364 17682
rect 55404 16652 55456 16658
rect 55404 16594 55456 16600
rect 56324 16652 56376 16658
rect 56324 16594 56376 16600
rect 55220 16584 55272 16590
rect 55220 16526 55272 16532
rect 55416 16250 55444 16594
rect 55496 16584 55548 16590
rect 55496 16526 55548 16532
rect 55404 16244 55456 16250
rect 55404 16186 55456 16192
rect 55036 16040 55088 16046
rect 55036 15982 55088 15988
rect 55508 15706 55536 16526
rect 55772 16108 55824 16114
rect 55772 16050 55824 16056
rect 55496 15700 55548 15706
rect 55496 15642 55548 15648
rect 54944 15632 54996 15638
rect 54944 15574 54996 15580
rect 55784 15502 55812 16050
rect 56336 15570 56364 16594
rect 56428 16114 56456 17818
rect 56704 17746 56732 18090
rect 56692 17740 56744 17746
rect 56692 17682 56744 17688
rect 57348 17610 57376 18702
rect 57428 18692 57480 18698
rect 57428 18634 57480 18640
rect 56784 17604 56836 17610
rect 56784 17546 56836 17552
rect 57336 17604 57388 17610
rect 57336 17546 57388 17552
rect 56692 17536 56744 17542
rect 56692 17478 56744 17484
rect 56704 16658 56732 17478
rect 56692 16652 56744 16658
rect 56692 16594 56744 16600
rect 56796 16454 56824 17546
rect 57242 17096 57298 17105
rect 57242 17031 57244 17040
rect 57296 17031 57298 17040
rect 57244 17002 57296 17008
rect 56600 16448 56652 16454
rect 56600 16390 56652 16396
rect 56784 16448 56836 16454
rect 56784 16390 56836 16396
rect 56416 16108 56468 16114
rect 56416 16050 56468 16056
rect 56612 15570 56640 16390
rect 57152 16108 57204 16114
rect 57152 16050 57204 16056
rect 57060 16040 57112 16046
rect 57058 16008 57060 16017
rect 57112 16008 57114 16017
rect 56692 15972 56744 15978
rect 57058 15943 57114 15952
rect 56692 15914 56744 15920
rect 56324 15564 56376 15570
rect 56324 15506 56376 15512
rect 56600 15564 56652 15570
rect 56600 15506 56652 15512
rect 55772 15496 55824 15502
rect 55772 15438 55824 15444
rect 56048 15088 56100 15094
rect 56048 15030 56100 15036
rect 54484 14408 54536 14414
rect 54484 14350 54536 14356
rect 54496 13938 54524 14350
rect 55588 14068 55640 14074
rect 55588 14010 55640 14016
rect 54484 13932 54536 13938
rect 54484 13874 54536 13880
rect 54116 12436 54168 12442
rect 54116 12378 54168 12384
rect 54392 12436 54444 12442
rect 54392 12378 54444 12384
rect 53932 11892 53984 11898
rect 53932 11834 53984 11840
rect 54128 11762 54156 12378
rect 54496 12306 54524 13874
rect 55600 13326 55628 14010
rect 56060 13802 56088 15030
rect 56704 14482 56732 15914
rect 56876 14952 56928 14958
rect 56876 14894 56928 14900
rect 56888 14618 56916 14894
rect 57164 14822 57192 16050
rect 57152 14816 57204 14822
rect 57152 14758 57204 14764
rect 57164 14618 57192 14758
rect 56876 14612 56928 14618
rect 56876 14554 56928 14560
rect 57152 14612 57204 14618
rect 57152 14554 57204 14560
rect 56692 14476 56744 14482
rect 56692 14418 56744 14424
rect 56140 14272 56192 14278
rect 56140 14214 56192 14220
rect 56152 13870 56180 14214
rect 57256 14074 57284 17002
rect 57440 16522 57468 18634
rect 57428 16516 57480 16522
rect 57428 16458 57480 16464
rect 57440 15586 57468 16458
rect 57348 15558 57468 15586
rect 57348 15434 57376 15558
rect 57336 15428 57388 15434
rect 57336 15370 57388 15376
rect 57348 14346 57376 15370
rect 57336 14340 57388 14346
rect 57336 14282 57388 14288
rect 57244 14068 57296 14074
rect 57244 14010 57296 14016
rect 56140 13864 56192 13870
rect 56140 13806 56192 13812
rect 56048 13796 56100 13802
rect 56048 13738 56100 13744
rect 55588 13320 55640 13326
rect 55588 13262 55640 13268
rect 55312 13184 55364 13190
rect 55312 13126 55364 13132
rect 55324 12918 55352 13126
rect 55312 12912 55364 12918
rect 55312 12854 55364 12860
rect 55600 12850 55628 13262
rect 55680 12980 55732 12986
rect 55680 12922 55732 12928
rect 55588 12844 55640 12850
rect 55588 12786 55640 12792
rect 55692 12782 55720 12922
rect 56060 12850 56088 13738
rect 56692 13728 56744 13734
rect 56692 13670 56744 13676
rect 56704 13394 56732 13670
rect 56692 13388 56744 13394
rect 56692 13330 56744 13336
rect 57348 13258 57376 14282
rect 57336 13252 57388 13258
rect 57336 13194 57388 13200
rect 56048 12844 56100 12850
rect 56048 12786 56100 12792
rect 57152 12844 57204 12850
rect 57152 12786 57204 12792
rect 55680 12776 55732 12782
rect 55680 12718 55732 12724
rect 54300 12300 54352 12306
rect 54300 12242 54352 12248
rect 54484 12300 54536 12306
rect 54484 12242 54536 12248
rect 53932 11756 53984 11762
rect 53852 11716 53932 11744
rect 53288 11698 53340 11704
rect 53932 11698 53984 11704
rect 54116 11756 54168 11762
rect 54116 11698 54168 11704
rect 51080 11688 51132 11694
rect 51080 11630 51132 11636
rect 52000 11688 52052 11694
rect 52000 11630 52052 11636
rect 53012 11688 53064 11694
rect 53012 11630 53064 11636
rect 53196 11688 53248 11694
rect 53196 11630 53248 11636
rect 51518 11452 51826 11461
rect 51518 11450 51524 11452
rect 51580 11450 51604 11452
rect 51660 11450 51684 11452
rect 51740 11450 51764 11452
rect 51820 11450 51826 11452
rect 51580 11398 51582 11450
rect 51762 11398 51764 11450
rect 51518 11396 51524 11398
rect 51580 11396 51604 11398
rect 51660 11396 51684 11398
rect 51740 11396 51764 11398
rect 51820 11396 51826 11398
rect 51518 11387 51826 11396
rect 52012 11082 52040 11630
rect 52644 11620 52696 11626
rect 52644 11562 52696 11568
rect 52092 11552 52144 11558
rect 52092 11494 52144 11500
rect 52104 11354 52132 11494
rect 52092 11348 52144 11354
rect 52092 11290 52144 11296
rect 52656 11150 52684 11562
rect 53104 11552 53156 11558
rect 53104 11494 53156 11500
rect 53116 11150 53144 11494
rect 53208 11354 53236 11630
rect 53196 11348 53248 11354
rect 53196 11290 53248 11296
rect 53300 11286 53328 11698
rect 53288 11280 53340 11286
rect 53288 11222 53340 11228
rect 53944 11150 53972 11698
rect 52644 11144 52696 11150
rect 52644 11086 52696 11092
rect 53104 11144 53156 11150
rect 53104 11086 53156 11092
rect 53932 11144 53984 11150
rect 53932 11086 53984 11092
rect 52000 11076 52052 11082
rect 52000 11018 52052 11024
rect 51908 11008 51960 11014
rect 51908 10950 51960 10956
rect 51920 10742 51948 10950
rect 52656 10810 52684 11086
rect 52644 10804 52696 10810
rect 52644 10746 52696 10752
rect 51908 10736 51960 10742
rect 51908 10678 51960 10684
rect 51356 10668 51408 10674
rect 51356 10610 51408 10616
rect 51080 10124 51132 10130
rect 51080 10066 51132 10072
rect 51092 9518 51120 10066
rect 51368 10062 51396 10610
rect 51448 10532 51500 10538
rect 51448 10474 51500 10480
rect 51356 10056 51408 10062
rect 51356 9998 51408 10004
rect 51460 9654 51488 10474
rect 51518 10364 51826 10373
rect 51518 10362 51524 10364
rect 51580 10362 51604 10364
rect 51660 10362 51684 10364
rect 51740 10362 51764 10364
rect 51820 10362 51826 10364
rect 51580 10310 51582 10362
rect 51762 10310 51764 10362
rect 51518 10308 51524 10310
rect 51580 10308 51604 10310
rect 51660 10308 51684 10310
rect 51740 10308 51764 10310
rect 51820 10308 51826 10310
rect 51518 10299 51826 10308
rect 51920 9994 51948 10678
rect 52368 10668 52420 10674
rect 52368 10610 52420 10616
rect 52380 10062 52408 10610
rect 53944 10266 53972 11086
rect 53932 10260 53984 10266
rect 53932 10202 53984 10208
rect 52368 10056 52420 10062
rect 52368 9998 52420 10004
rect 52644 10056 52696 10062
rect 52644 9998 52696 10004
rect 51908 9988 51960 9994
rect 51908 9930 51960 9936
rect 52656 9654 52684 9998
rect 51448 9648 51500 9654
rect 51448 9590 51500 9596
rect 52644 9648 52696 9654
rect 52644 9590 52696 9596
rect 54312 9586 54340 12242
rect 55692 12238 55720 12718
rect 56600 12708 56652 12714
rect 56600 12650 56652 12656
rect 55680 12232 55732 12238
rect 55680 12174 55732 12180
rect 55312 12096 55364 12102
rect 55312 12038 55364 12044
rect 55324 11762 55352 12038
rect 54944 11756 54996 11762
rect 54944 11698 54996 11704
rect 55312 11756 55364 11762
rect 55312 11698 55364 11704
rect 54956 11354 54984 11698
rect 56140 11688 56192 11694
rect 56140 11630 56192 11636
rect 54944 11348 54996 11354
rect 54944 11290 54996 11296
rect 56152 11218 56180 11630
rect 56140 11212 56192 11218
rect 56140 11154 56192 11160
rect 56612 11082 56640 12650
rect 56784 12164 56836 12170
rect 56784 12106 56836 12112
rect 56796 11898 56824 12106
rect 56784 11892 56836 11898
rect 56784 11834 56836 11840
rect 57164 11354 57192 12786
rect 57152 11348 57204 11354
rect 57152 11290 57204 11296
rect 56600 11076 56652 11082
rect 56600 11018 56652 11024
rect 56048 10668 56100 10674
rect 56048 10610 56100 10616
rect 54576 10532 54628 10538
rect 54576 10474 54628 10480
rect 54588 9654 54616 10474
rect 55404 10192 55456 10198
rect 55404 10134 55456 10140
rect 55128 10124 55180 10130
rect 55128 10066 55180 10072
rect 54576 9648 54628 9654
rect 54576 9590 54628 9596
rect 54300 9580 54352 9586
rect 54300 9522 54352 9528
rect 51080 9512 51132 9518
rect 51080 9454 51132 9460
rect 51518 9276 51826 9285
rect 51518 9274 51524 9276
rect 51580 9274 51604 9276
rect 51660 9274 51684 9276
rect 51740 9274 51764 9276
rect 51820 9274 51826 9276
rect 51580 9222 51582 9274
rect 51762 9222 51764 9274
rect 51518 9220 51524 9222
rect 51580 9220 51604 9222
rect 51660 9220 51684 9222
rect 51740 9220 51764 9222
rect 51820 9220 51826 9222
rect 51518 9211 51826 9220
rect 55140 9178 55168 10066
rect 55416 9625 55444 10134
rect 55402 9616 55458 9625
rect 55402 9551 55458 9560
rect 50988 9172 51040 9178
rect 50988 9114 51040 9120
rect 55128 9172 55180 9178
rect 55128 9114 55180 9120
rect 55416 8634 55444 9551
rect 56060 9518 56088 10610
rect 56612 10130 56640 11018
rect 56600 10124 56652 10130
rect 56600 10066 56652 10072
rect 57336 10124 57388 10130
rect 57336 10066 57388 10072
rect 56612 9654 56640 10066
rect 56600 9648 56652 9654
rect 56600 9590 56652 9596
rect 56048 9512 56100 9518
rect 56048 9454 56100 9460
rect 55586 8936 55642 8945
rect 56612 8906 56640 9590
rect 57348 9042 57376 10066
rect 57532 9994 57560 33254
rect 57808 33114 57836 33458
rect 58070 33416 58126 33425
rect 58070 33351 58072 33360
rect 58124 33351 58126 33360
rect 58072 33322 58124 33328
rect 57796 33108 57848 33114
rect 57796 33050 57848 33056
rect 58072 28076 58124 28082
rect 58072 28018 58124 28024
rect 58084 27985 58112 28018
rect 58070 27976 58126 27985
rect 57704 27940 57756 27946
rect 58070 27911 58126 27920
rect 57704 27882 57756 27888
rect 57716 12434 57744 27882
rect 58084 27674 58112 27911
rect 58072 27668 58124 27674
rect 58072 27610 58124 27616
rect 57888 23520 57940 23526
rect 57888 23462 57940 23468
rect 57900 23225 57928 23462
rect 57886 23216 57942 23225
rect 57886 23151 57942 23160
rect 57888 18284 57940 18290
rect 57888 18226 57940 18232
rect 57796 18080 57848 18086
rect 57796 18022 57848 18028
rect 57808 17785 57836 18022
rect 57794 17776 57850 17785
rect 57794 17711 57850 17720
rect 57900 17338 57928 18226
rect 57888 17332 57940 17338
rect 57888 17274 57940 17280
rect 57980 13932 58032 13938
rect 57980 13874 58032 13880
rect 57888 13728 57940 13734
rect 57888 13670 57940 13676
rect 57624 12406 57744 12434
rect 57624 11121 57652 12406
rect 57796 11552 57848 11558
rect 57796 11494 57848 11500
rect 57808 11218 57836 11494
rect 57796 11212 57848 11218
rect 57796 11154 57848 11160
rect 57610 11112 57666 11121
rect 57610 11047 57666 11056
rect 57520 9988 57572 9994
rect 57520 9930 57572 9936
rect 57532 9722 57560 9930
rect 57520 9716 57572 9722
rect 57520 9658 57572 9664
rect 57336 9036 57388 9042
rect 57336 8978 57388 8984
rect 55586 8871 55642 8880
rect 56600 8900 56652 8906
rect 55600 8838 55628 8871
rect 56600 8842 56652 8848
rect 55588 8832 55640 8838
rect 55588 8774 55640 8780
rect 57796 8832 57848 8838
rect 57796 8774 57848 8780
rect 55404 8628 55456 8634
rect 55404 8570 55456 8576
rect 51518 8188 51826 8197
rect 51518 8186 51524 8188
rect 51580 8186 51604 8188
rect 51660 8186 51684 8188
rect 51740 8186 51764 8188
rect 51820 8186 51826 8188
rect 51580 8134 51582 8186
rect 51762 8134 51764 8186
rect 51518 8132 51524 8134
rect 51580 8132 51604 8134
rect 51660 8132 51684 8134
rect 51740 8132 51764 8134
rect 51820 8132 51826 8134
rect 51518 8123 51826 8132
rect 57808 8022 57836 8774
rect 57796 8016 57848 8022
rect 57796 7958 57848 7964
rect 51518 7100 51826 7109
rect 51518 7098 51524 7100
rect 51580 7098 51604 7100
rect 51660 7098 51684 7100
rect 51740 7098 51764 7100
rect 51820 7098 51826 7100
rect 51580 7046 51582 7098
rect 51762 7046 51764 7098
rect 51518 7044 51524 7046
rect 51580 7044 51604 7046
rect 51660 7044 51684 7046
rect 51740 7044 51764 7046
rect 51820 7044 51826 7046
rect 51518 7035 51826 7044
rect 51518 6012 51826 6021
rect 51518 6010 51524 6012
rect 51580 6010 51604 6012
rect 51660 6010 51684 6012
rect 51740 6010 51764 6012
rect 51820 6010 51826 6012
rect 51580 5958 51582 6010
rect 51762 5958 51764 6010
rect 51518 5956 51524 5958
rect 51580 5956 51604 5958
rect 51660 5956 51684 5958
rect 51740 5956 51764 5958
rect 51820 5956 51826 5958
rect 51518 5947 51826 5956
rect 51518 4924 51826 4933
rect 51518 4922 51524 4924
rect 51580 4922 51604 4924
rect 51660 4922 51684 4924
rect 51740 4922 51764 4924
rect 51820 4922 51826 4924
rect 51580 4870 51582 4922
rect 51762 4870 51764 4922
rect 51518 4868 51524 4870
rect 51580 4868 51604 4870
rect 51660 4868 51684 4870
rect 51740 4868 51764 4870
rect 51820 4868 51826 4870
rect 51518 4859 51826 4868
rect 48688 4140 48740 4146
rect 48688 4082 48740 4088
rect 48700 3738 48728 4082
rect 48872 3936 48924 3942
rect 48872 3878 48924 3884
rect 48688 3732 48740 3738
rect 48688 3674 48740 3680
rect 48884 3058 48912 3878
rect 51518 3836 51826 3845
rect 51518 3834 51524 3836
rect 51580 3834 51604 3836
rect 51660 3834 51684 3836
rect 51740 3834 51764 3836
rect 51820 3834 51826 3836
rect 51580 3782 51582 3834
rect 51762 3782 51764 3834
rect 51518 3780 51524 3782
rect 51580 3780 51604 3782
rect 51660 3780 51684 3782
rect 51740 3780 51764 3782
rect 51820 3780 51826 3782
rect 51518 3771 51826 3780
rect 48872 3052 48924 3058
rect 48872 2994 48924 3000
rect 53104 2916 53156 2922
rect 53104 2858 53156 2864
rect 52828 2848 52880 2854
rect 52828 2790 52880 2796
rect 51518 2748 51826 2757
rect 51518 2746 51524 2748
rect 51580 2746 51604 2748
rect 51660 2746 51684 2748
rect 51740 2746 51764 2748
rect 51820 2746 51826 2748
rect 51580 2694 51582 2746
rect 51762 2694 51764 2746
rect 51518 2692 51524 2694
rect 51580 2692 51604 2694
rect 51660 2692 51684 2694
rect 51740 2692 51764 2694
rect 51820 2692 51826 2694
rect 51518 2683 51826 2692
rect 43168 2440 43220 2446
rect 43168 2382 43220 2388
rect 48412 2440 48464 2446
rect 48412 2382 48464 2388
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 41420 2372 41472 2378
rect 41420 2314 41472 2320
rect 9692 800 9720 2314
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 29000 2304 29052 2310
rect 29000 2246 29052 2252
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 14200 800 14228 2246
rect 15398 2204 15706 2213
rect 15398 2202 15404 2204
rect 15460 2202 15484 2204
rect 15540 2202 15564 2204
rect 15620 2202 15644 2204
rect 15700 2202 15706 2204
rect 15460 2150 15462 2202
rect 15642 2150 15644 2202
rect 15398 2148 15404 2150
rect 15460 2148 15484 2150
rect 15540 2148 15564 2150
rect 15620 2148 15644 2150
rect 15700 2148 15706 2150
rect 15398 2139 15706 2148
rect 19352 800 19380 2246
rect 23860 800 23888 2246
rect 29012 800 29040 2246
rect 29846 2204 30154 2213
rect 29846 2202 29852 2204
rect 29908 2202 29932 2204
rect 29988 2202 30012 2204
rect 30068 2202 30092 2204
rect 30148 2202 30154 2204
rect 29908 2150 29910 2202
rect 30090 2150 30092 2202
rect 29846 2148 29852 2150
rect 29908 2148 29932 2150
rect 29988 2148 30012 2150
rect 30068 2148 30092 2150
rect 30148 2148 30154 2150
rect 29846 2139 30154 2148
rect 33520 800 33548 2246
rect 38672 800 38700 2246
rect 43180 800 43208 2382
rect 52840 2378 52868 2790
rect 53116 2582 53144 2858
rect 53104 2576 53156 2582
rect 53104 2518 53156 2524
rect 57900 2446 57928 13670
rect 57992 13530 58020 13874
rect 57980 13524 58032 13530
rect 57980 13466 58032 13472
rect 58070 13016 58126 13025
rect 58070 12951 58072 12960
rect 58124 12951 58126 12960
rect 58072 12922 58124 12928
rect 58072 7812 58124 7818
rect 58072 7754 58124 7760
rect 58084 7585 58112 7754
rect 58070 7576 58126 7585
rect 58070 7511 58126 7520
rect 58072 2848 58124 2854
rect 58070 2816 58072 2825
rect 58124 2816 58126 2825
rect 58070 2751 58126 2760
rect 57888 2440 57940 2446
rect 57888 2382 57940 2388
rect 52828 2372 52880 2378
rect 52828 2314 52880 2320
rect 48320 2304 48372 2310
rect 48320 2246 48372 2252
rect 44294 2204 44602 2213
rect 44294 2202 44300 2204
rect 44356 2202 44380 2204
rect 44436 2202 44460 2204
rect 44516 2202 44540 2204
rect 44596 2202 44602 2204
rect 44356 2150 44358 2202
rect 44538 2150 44540 2202
rect 44294 2148 44300 2150
rect 44356 2148 44380 2150
rect 44436 2148 44460 2150
rect 44516 2148 44540 2150
rect 44596 2148 44602 2150
rect 44294 2139 44602 2148
rect 48332 800 48360 2246
rect 52840 800 52868 2314
rect 57980 2304 58032 2310
rect 57980 2246 58032 2252
rect 57992 800 58020 2246
rect 18 0 74 800
rect 4526 0 4582 800
rect 9678 0 9734 800
rect 14186 0 14242 800
rect 19338 0 19394 800
rect 23846 0 23902 800
rect 28998 0 29054 800
rect 33506 0 33562 800
rect 38658 0 38714 800
rect 43166 0 43222 800
rect 48318 0 48374 800
rect 52826 0 52882 800
rect 57978 0 58034 800
<< via2 >>
rect 1490 35400 1546 35456
rect 15404 33754 15460 33756
rect 15484 33754 15540 33756
rect 15564 33754 15620 33756
rect 15644 33754 15700 33756
rect 15404 33702 15450 33754
rect 15450 33702 15460 33754
rect 15484 33702 15514 33754
rect 15514 33702 15526 33754
rect 15526 33702 15540 33754
rect 15564 33702 15578 33754
rect 15578 33702 15590 33754
rect 15590 33702 15620 33754
rect 15644 33702 15654 33754
rect 15654 33702 15700 33754
rect 15404 33700 15460 33702
rect 15484 33700 15540 33702
rect 15564 33700 15620 33702
rect 15644 33700 15700 33702
rect 29852 33754 29908 33756
rect 29932 33754 29988 33756
rect 30012 33754 30068 33756
rect 30092 33754 30148 33756
rect 29852 33702 29898 33754
rect 29898 33702 29908 33754
rect 29932 33702 29962 33754
rect 29962 33702 29974 33754
rect 29974 33702 29988 33754
rect 30012 33702 30026 33754
rect 30026 33702 30038 33754
rect 30038 33702 30068 33754
rect 30092 33702 30102 33754
rect 30102 33702 30148 33754
rect 29852 33700 29908 33702
rect 29932 33700 29988 33702
rect 30012 33700 30068 33702
rect 30092 33700 30148 33702
rect 44300 33754 44356 33756
rect 44380 33754 44436 33756
rect 44460 33754 44516 33756
rect 44540 33754 44596 33756
rect 44300 33702 44346 33754
rect 44346 33702 44356 33754
rect 44380 33702 44410 33754
rect 44410 33702 44422 33754
rect 44422 33702 44436 33754
rect 44460 33702 44474 33754
rect 44474 33702 44486 33754
rect 44486 33702 44516 33754
rect 44540 33702 44550 33754
rect 44550 33702 44596 33754
rect 44300 33700 44356 33702
rect 44380 33700 44436 33702
rect 44460 33700 44516 33702
rect 44540 33700 44596 33702
rect 1490 30640 1546 30696
rect 1490 25200 1546 25256
rect 2410 24792 2466 24848
rect 4250 27920 4306 27976
rect 2042 23160 2098 23216
rect 2962 20440 3018 20496
rect 3974 18264 4030 18320
rect 4066 18128 4122 18184
rect 5814 23568 5870 23624
rect 4894 23024 4950 23080
rect 4618 16224 4674 16280
rect 4894 16088 4950 16144
rect 5722 15408 5778 15464
rect 5446 14864 5502 14920
rect 3790 14320 3846 14376
rect 7378 22616 7434 22672
rect 6274 16496 6330 16552
rect 6458 15972 6514 16008
rect 6458 15952 6460 15972
rect 6460 15952 6512 15972
rect 6512 15952 6514 15972
rect 8180 33210 8236 33212
rect 8260 33210 8316 33212
rect 8340 33210 8396 33212
rect 8420 33210 8476 33212
rect 8180 33158 8226 33210
rect 8226 33158 8236 33210
rect 8260 33158 8290 33210
rect 8290 33158 8302 33210
rect 8302 33158 8316 33210
rect 8340 33158 8354 33210
rect 8354 33158 8366 33210
rect 8366 33158 8396 33210
rect 8420 33158 8430 33210
rect 8430 33158 8476 33210
rect 8180 33156 8236 33158
rect 8260 33156 8316 33158
rect 8340 33156 8396 33158
rect 8420 33156 8476 33158
rect 15404 32666 15460 32668
rect 15484 32666 15540 32668
rect 15564 32666 15620 32668
rect 15644 32666 15700 32668
rect 15404 32614 15450 32666
rect 15450 32614 15460 32666
rect 15484 32614 15514 32666
rect 15514 32614 15526 32666
rect 15526 32614 15540 32666
rect 15564 32614 15578 32666
rect 15578 32614 15590 32666
rect 15590 32614 15620 32666
rect 15644 32614 15654 32666
rect 15654 32614 15700 32666
rect 15404 32612 15460 32614
rect 15484 32612 15540 32614
rect 15564 32612 15620 32614
rect 15644 32612 15700 32614
rect 8180 32122 8236 32124
rect 8260 32122 8316 32124
rect 8340 32122 8396 32124
rect 8420 32122 8476 32124
rect 8180 32070 8226 32122
rect 8226 32070 8236 32122
rect 8260 32070 8290 32122
rect 8290 32070 8302 32122
rect 8302 32070 8316 32122
rect 8340 32070 8354 32122
rect 8354 32070 8366 32122
rect 8366 32070 8396 32122
rect 8420 32070 8430 32122
rect 8430 32070 8476 32122
rect 8180 32068 8236 32070
rect 8260 32068 8316 32070
rect 8340 32068 8396 32070
rect 8420 32068 8476 32070
rect 8180 31034 8236 31036
rect 8260 31034 8316 31036
rect 8340 31034 8396 31036
rect 8420 31034 8476 31036
rect 8180 30982 8226 31034
rect 8226 30982 8236 31034
rect 8260 30982 8290 31034
rect 8290 30982 8302 31034
rect 8302 30982 8316 31034
rect 8340 30982 8354 31034
rect 8354 30982 8366 31034
rect 8366 30982 8396 31034
rect 8420 30982 8430 31034
rect 8430 30982 8476 31034
rect 8180 30980 8236 30982
rect 8260 30980 8316 30982
rect 8340 30980 8396 30982
rect 8420 30980 8476 30982
rect 8180 29946 8236 29948
rect 8260 29946 8316 29948
rect 8340 29946 8396 29948
rect 8420 29946 8476 29948
rect 8180 29894 8226 29946
rect 8226 29894 8236 29946
rect 8260 29894 8290 29946
rect 8290 29894 8302 29946
rect 8302 29894 8316 29946
rect 8340 29894 8354 29946
rect 8354 29894 8366 29946
rect 8366 29894 8396 29946
rect 8420 29894 8430 29946
rect 8430 29894 8476 29946
rect 8180 29892 8236 29894
rect 8260 29892 8316 29894
rect 8340 29892 8396 29894
rect 8420 29892 8476 29894
rect 8180 28858 8236 28860
rect 8260 28858 8316 28860
rect 8340 28858 8396 28860
rect 8420 28858 8476 28860
rect 8180 28806 8226 28858
rect 8226 28806 8236 28858
rect 8260 28806 8290 28858
rect 8290 28806 8302 28858
rect 8302 28806 8316 28858
rect 8340 28806 8354 28858
rect 8354 28806 8366 28858
rect 8366 28806 8396 28858
rect 8420 28806 8430 28858
rect 8430 28806 8476 28858
rect 8180 28804 8236 28806
rect 8260 28804 8316 28806
rect 8340 28804 8396 28806
rect 8420 28804 8476 28806
rect 8180 27770 8236 27772
rect 8260 27770 8316 27772
rect 8340 27770 8396 27772
rect 8420 27770 8476 27772
rect 8180 27718 8226 27770
rect 8226 27718 8236 27770
rect 8260 27718 8290 27770
rect 8290 27718 8302 27770
rect 8302 27718 8316 27770
rect 8340 27718 8354 27770
rect 8354 27718 8366 27770
rect 8366 27718 8396 27770
rect 8420 27718 8430 27770
rect 8430 27718 8476 27770
rect 8180 27716 8236 27718
rect 8260 27716 8316 27718
rect 8340 27716 8396 27718
rect 8420 27716 8476 27718
rect 8180 26682 8236 26684
rect 8260 26682 8316 26684
rect 8340 26682 8396 26684
rect 8420 26682 8476 26684
rect 8180 26630 8226 26682
rect 8226 26630 8236 26682
rect 8260 26630 8290 26682
rect 8290 26630 8302 26682
rect 8302 26630 8316 26682
rect 8340 26630 8354 26682
rect 8354 26630 8366 26682
rect 8366 26630 8396 26682
rect 8420 26630 8430 26682
rect 8430 26630 8476 26682
rect 8180 26628 8236 26630
rect 8260 26628 8316 26630
rect 8340 26628 8396 26630
rect 8420 26628 8476 26630
rect 8180 25594 8236 25596
rect 8260 25594 8316 25596
rect 8340 25594 8396 25596
rect 8420 25594 8476 25596
rect 8180 25542 8226 25594
rect 8226 25542 8236 25594
rect 8260 25542 8290 25594
rect 8290 25542 8302 25594
rect 8302 25542 8316 25594
rect 8340 25542 8354 25594
rect 8354 25542 8366 25594
rect 8366 25542 8396 25594
rect 8420 25542 8430 25594
rect 8430 25542 8476 25594
rect 8180 25540 8236 25542
rect 8260 25540 8316 25542
rect 8340 25540 8396 25542
rect 8420 25540 8476 25542
rect 8180 24506 8236 24508
rect 8260 24506 8316 24508
rect 8340 24506 8396 24508
rect 8420 24506 8476 24508
rect 8180 24454 8226 24506
rect 8226 24454 8236 24506
rect 8260 24454 8290 24506
rect 8290 24454 8302 24506
rect 8302 24454 8316 24506
rect 8340 24454 8354 24506
rect 8354 24454 8366 24506
rect 8366 24454 8396 24506
rect 8420 24454 8430 24506
rect 8430 24454 8476 24506
rect 8180 24452 8236 24454
rect 8260 24452 8316 24454
rect 8340 24452 8396 24454
rect 8420 24452 8476 24454
rect 8114 24268 8170 24304
rect 8114 24248 8116 24268
rect 8116 24248 8168 24268
rect 8168 24248 8170 24268
rect 8180 23418 8236 23420
rect 8260 23418 8316 23420
rect 8340 23418 8396 23420
rect 8420 23418 8476 23420
rect 8180 23366 8226 23418
rect 8226 23366 8236 23418
rect 8260 23366 8290 23418
rect 8290 23366 8302 23418
rect 8302 23366 8316 23418
rect 8340 23366 8354 23418
rect 8354 23366 8366 23418
rect 8366 23366 8396 23418
rect 8420 23366 8430 23418
rect 8430 23366 8476 23418
rect 8180 23364 8236 23366
rect 8260 23364 8316 23366
rect 8340 23364 8396 23366
rect 8420 23364 8476 23366
rect 8180 22330 8236 22332
rect 8260 22330 8316 22332
rect 8340 22330 8396 22332
rect 8420 22330 8476 22332
rect 8180 22278 8226 22330
rect 8226 22278 8236 22330
rect 8260 22278 8290 22330
rect 8290 22278 8302 22330
rect 8302 22278 8316 22330
rect 8340 22278 8354 22330
rect 8354 22278 8366 22330
rect 8366 22278 8396 22330
rect 8420 22278 8430 22330
rect 8430 22278 8476 22330
rect 8180 22276 8236 22278
rect 8260 22276 8316 22278
rect 8340 22276 8396 22278
rect 8420 22276 8476 22278
rect 8180 21242 8236 21244
rect 8260 21242 8316 21244
rect 8340 21242 8396 21244
rect 8420 21242 8476 21244
rect 8180 21190 8226 21242
rect 8226 21190 8236 21242
rect 8260 21190 8290 21242
rect 8290 21190 8302 21242
rect 8302 21190 8316 21242
rect 8340 21190 8354 21242
rect 8354 21190 8366 21242
rect 8366 21190 8396 21242
rect 8420 21190 8430 21242
rect 8430 21190 8476 21242
rect 8180 21188 8236 21190
rect 8260 21188 8316 21190
rect 8340 21188 8396 21190
rect 8420 21188 8476 21190
rect 8180 20154 8236 20156
rect 8260 20154 8316 20156
rect 8340 20154 8396 20156
rect 8420 20154 8476 20156
rect 8180 20102 8226 20154
rect 8226 20102 8236 20154
rect 8260 20102 8290 20154
rect 8290 20102 8302 20154
rect 8302 20102 8316 20154
rect 8340 20102 8354 20154
rect 8354 20102 8366 20154
rect 8366 20102 8396 20154
rect 8420 20102 8430 20154
rect 8430 20102 8476 20154
rect 8180 20100 8236 20102
rect 8260 20100 8316 20102
rect 8340 20100 8396 20102
rect 8420 20100 8476 20102
rect 8180 19066 8236 19068
rect 8260 19066 8316 19068
rect 8340 19066 8396 19068
rect 8420 19066 8476 19068
rect 8180 19014 8226 19066
rect 8226 19014 8236 19066
rect 8260 19014 8290 19066
rect 8290 19014 8302 19066
rect 8302 19014 8316 19066
rect 8340 19014 8354 19066
rect 8354 19014 8366 19066
rect 8366 19014 8396 19066
rect 8420 19014 8430 19066
rect 8430 19014 8476 19066
rect 8180 19012 8236 19014
rect 8260 19012 8316 19014
rect 8340 19012 8396 19014
rect 8420 19012 8476 19014
rect 8180 17978 8236 17980
rect 8260 17978 8316 17980
rect 8340 17978 8396 17980
rect 8420 17978 8476 17980
rect 8180 17926 8226 17978
rect 8226 17926 8236 17978
rect 8260 17926 8290 17978
rect 8290 17926 8302 17978
rect 8302 17926 8316 17978
rect 8340 17926 8354 17978
rect 8354 17926 8366 17978
rect 8366 17926 8396 17978
rect 8420 17926 8430 17978
rect 8430 17926 8476 17978
rect 8180 17924 8236 17926
rect 8260 17924 8316 17926
rect 8340 17924 8396 17926
rect 8420 17924 8476 17926
rect 8180 16890 8236 16892
rect 8260 16890 8316 16892
rect 8340 16890 8396 16892
rect 8420 16890 8476 16892
rect 8180 16838 8226 16890
rect 8226 16838 8236 16890
rect 8260 16838 8290 16890
rect 8290 16838 8302 16890
rect 8302 16838 8316 16890
rect 8340 16838 8354 16890
rect 8354 16838 8366 16890
rect 8366 16838 8396 16890
rect 8420 16838 8430 16890
rect 8430 16838 8476 16890
rect 8180 16836 8236 16838
rect 8260 16836 8316 16838
rect 8340 16836 8396 16838
rect 8420 16836 8476 16838
rect 6458 13232 6514 13288
rect 5814 12280 5870 12336
rect 1582 10260 1638 10296
rect 1582 10240 1584 10260
rect 1584 10240 1636 10260
rect 1636 10240 1638 10260
rect 1490 4800 1546 4856
rect 8180 15802 8236 15804
rect 8260 15802 8316 15804
rect 8340 15802 8396 15804
rect 8420 15802 8476 15804
rect 8180 15750 8226 15802
rect 8226 15750 8236 15802
rect 8260 15750 8290 15802
rect 8290 15750 8302 15802
rect 8302 15750 8316 15802
rect 8340 15750 8354 15802
rect 8354 15750 8366 15802
rect 8366 15750 8396 15802
rect 8420 15750 8430 15802
rect 8430 15750 8476 15802
rect 8180 15748 8236 15750
rect 8260 15748 8316 15750
rect 8340 15748 8396 15750
rect 8420 15748 8476 15750
rect 8298 15564 8354 15600
rect 8298 15544 8300 15564
rect 8300 15544 8352 15564
rect 8352 15544 8354 15564
rect 15404 31578 15460 31580
rect 15484 31578 15540 31580
rect 15564 31578 15620 31580
rect 15644 31578 15700 31580
rect 15404 31526 15450 31578
rect 15450 31526 15460 31578
rect 15484 31526 15514 31578
rect 15514 31526 15526 31578
rect 15526 31526 15540 31578
rect 15564 31526 15578 31578
rect 15578 31526 15590 31578
rect 15590 31526 15620 31578
rect 15644 31526 15654 31578
rect 15654 31526 15700 31578
rect 15404 31524 15460 31526
rect 15484 31524 15540 31526
rect 15564 31524 15620 31526
rect 15644 31524 15700 31526
rect 15404 30490 15460 30492
rect 15484 30490 15540 30492
rect 15564 30490 15620 30492
rect 15644 30490 15700 30492
rect 15404 30438 15450 30490
rect 15450 30438 15460 30490
rect 15484 30438 15514 30490
rect 15514 30438 15526 30490
rect 15526 30438 15540 30490
rect 15564 30438 15578 30490
rect 15578 30438 15590 30490
rect 15590 30438 15620 30490
rect 15644 30438 15654 30490
rect 15654 30438 15700 30490
rect 15404 30436 15460 30438
rect 15484 30436 15540 30438
rect 15564 30436 15620 30438
rect 15644 30436 15700 30438
rect 9034 27920 9090 27976
rect 15404 29402 15460 29404
rect 15484 29402 15540 29404
rect 15564 29402 15620 29404
rect 15644 29402 15700 29404
rect 15404 29350 15450 29402
rect 15450 29350 15460 29402
rect 15484 29350 15514 29402
rect 15514 29350 15526 29402
rect 15526 29350 15540 29402
rect 15564 29350 15578 29402
rect 15578 29350 15590 29402
rect 15590 29350 15620 29402
rect 15644 29350 15654 29402
rect 15654 29350 15700 29402
rect 15404 29348 15460 29350
rect 15484 29348 15540 29350
rect 15564 29348 15620 29350
rect 15644 29348 15700 29350
rect 15404 28314 15460 28316
rect 15484 28314 15540 28316
rect 15564 28314 15620 28316
rect 15644 28314 15700 28316
rect 15404 28262 15450 28314
rect 15450 28262 15460 28314
rect 15484 28262 15514 28314
rect 15514 28262 15526 28314
rect 15526 28262 15540 28314
rect 15564 28262 15578 28314
rect 15578 28262 15590 28314
rect 15590 28262 15620 28314
rect 15644 28262 15654 28314
rect 15654 28262 15700 28314
rect 15404 28260 15460 28262
rect 15484 28260 15540 28262
rect 15564 28260 15620 28262
rect 15644 28260 15700 28262
rect 15404 27226 15460 27228
rect 15484 27226 15540 27228
rect 15564 27226 15620 27228
rect 15644 27226 15700 27228
rect 15404 27174 15450 27226
rect 15450 27174 15460 27226
rect 15484 27174 15514 27226
rect 15514 27174 15526 27226
rect 15526 27174 15540 27226
rect 15564 27174 15578 27226
rect 15578 27174 15590 27226
rect 15590 27174 15620 27226
rect 15644 27174 15654 27226
rect 15654 27174 15700 27226
rect 15404 27172 15460 27174
rect 15484 27172 15540 27174
rect 15564 27172 15620 27174
rect 15644 27172 15700 27174
rect 8180 14714 8236 14716
rect 8260 14714 8316 14716
rect 8340 14714 8396 14716
rect 8420 14714 8476 14716
rect 8180 14662 8226 14714
rect 8226 14662 8236 14714
rect 8260 14662 8290 14714
rect 8290 14662 8302 14714
rect 8302 14662 8316 14714
rect 8340 14662 8354 14714
rect 8354 14662 8366 14714
rect 8366 14662 8396 14714
rect 8420 14662 8430 14714
rect 8430 14662 8476 14714
rect 8180 14660 8236 14662
rect 8260 14660 8316 14662
rect 8340 14660 8396 14662
rect 8420 14660 8476 14662
rect 8298 14492 8300 14512
rect 8300 14492 8352 14512
rect 8352 14492 8354 14512
rect 8298 14456 8354 14492
rect 9310 17720 9366 17776
rect 9126 16224 9182 16280
rect 8758 13932 8814 13968
rect 8758 13912 8760 13932
rect 8760 13912 8812 13932
rect 8812 13912 8814 13932
rect 8180 13626 8236 13628
rect 8260 13626 8316 13628
rect 8340 13626 8396 13628
rect 8420 13626 8476 13628
rect 8180 13574 8226 13626
rect 8226 13574 8236 13626
rect 8260 13574 8290 13626
rect 8290 13574 8302 13626
rect 8302 13574 8316 13626
rect 8340 13574 8354 13626
rect 8354 13574 8366 13626
rect 8366 13574 8396 13626
rect 8420 13574 8430 13626
rect 8430 13574 8476 13626
rect 8180 13572 8236 13574
rect 8260 13572 8316 13574
rect 8340 13572 8396 13574
rect 8420 13572 8476 13574
rect 8180 12538 8236 12540
rect 8260 12538 8316 12540
rect 8340 12538 8396 12540
rect 8420 12538 8476 12540
rect 8180 12486 8226 12538
rect 8226 12486 8236 12538
rect 8260 12486 8290 12538
rect 8290 12486 8302 12538
rect 8302 12486 8316 12538
rect 8340 12486 8354 12538
rect 8354 12486 8366 12538
rect 8366 12486 8396 12538
rect 8420 12486 8430 12538
rect 8430 12486 8476 12538
rect 8180 12484 8236 12486
rect 8260 12484 8316 12486
rect 8340 12484 8396 12486
rect 8420 12484 8476 12486
rect 12622 25356 12678 25392
rect 12622 25336 12624 25356
rect 12624 25336 12676 25356
rect 12676 25336 12678 25356
rect 13634 24112 13690 24168
rect 12070 17040 12126 17096
rect 8180 11450 8236 11452
rect 8260 11450 8316 11452
rect 8340 11450 8396 11452
rect 8420 11450 8476 11452
rect 8180 11398 8226 11450
rect 8226 11398 8236 11450
rect 8260 11398 8290 11450
rect 8290 11398 8302 11450
rect 8302 11398 8316 11450
rect 8340 11398 8354 11450
rect 8354 11398 8366 11450
rect 8366 11398 8396 11450
rect 8420 11398 8430 11450
rect 8430 11398 8476 11450
rect 8180 11396 8236 11398
rect 8260 11396 8316 11398
rect 8340 11396 8396 11398
rect 8420 11396 8476 11398
rect 12622 12844 12678 12880
rect 12622 12824 12624 12844
rect 12624 12824 12676 12844
rect 12676 12824 12678 12844
rect 13542 11736 13598 11792
rect 8180 10362 8236 10364
rect 8260 10362 8316 10364
rect 8340 10362 8396 10364
rect 8420 10362 8476 10364
rect 8180 10310 8226 10362
rect 8226 10310 8236 10362
rect 8260 10310 8290 10362
rect 8290 10310 8302 10362
rect 8302 10310 8316 10362
rect 8340 10310 8354 10362
rect 8354 10310 8366 10362
rect 8366 10310 8396 10362
rect 8420 10310 8430 10362
rect 8430 10310 8476 10362
rect 8180 10308 8236 10310
rect 8260 10308 8316 10310
rect 8340 10308 8396 10310
rect 8420 10308 8476 10310
rect 8180 9274 8236 9276
rect 8260 9274 8316 9276
rect 8340 9274 8396 9276
rect 8420 9274 8476 9276
rect 8180 9222 8226 9274
rect 8226 9222 8236 9274
rect 8260 9222 8290 9274
rect 8290 9222 8302 9274
rect 8302 9222 8316 9274
rect 8340 9222 8354 9274
rect 8354 9222 8366 9274
rect 8366 9222 8396 9274
rect 8420 9222 8430 9274
rect 8430 9222 8476 9274
rect 8180 9220 8236 9222
rect 8260 9220 8316 9222
rect 8340 9220 8396 9222
rect 8420 9220 8476 9222
rect 8180 8186 8236 8188
rect 8260 8186 8316 8188
rect 8340 8186 8396 8188
rect 8420 8186 8476 8188
rect 8180 8134 8226 8186
rect 8226 8134 8236 8186
rect 8260 8134 8290 8186
rect 8290 8134 8302 8186
rect 8302 8134 8316 8186
rect 8340 8134 8354 8186
rect 8354 8134 8366 8186
rect 8366 8134 8396 8186
rect 8420 8134 8430 8186
rect 8430 8134 8476 8186
rect 8180 8132 8236 8134
rect 8260 8132 8316 8134
rect 8340 8132 8396 8134
rect 8420 8132 8476 8134
rect 8180 7098 8236 7100
rect 8260 7098 8316 7100
rect 8340 7098 8396 7100
rect 8420 7098 8476 7100
rect 8180 7046 8226 7098
rect 8226 7046 8236 7098
rect 8260 7046 8290 7098
rect 8290 7046 8302 7098
rect 8302 7046 8316 7098
rect 8340 7046 8354 7098
rect 8354 7046 8366 7098
rect 8366 7046 8396 7098
rect 8420 7046 8430 7098
rect 8430 7046 8476 7098
rect 8180 7044 8236 7046
rect 8260 7044 8316 7046
rect 8340 7044 8396 7046
rect 8420 7044 8476 7046
rect 8180 6010 8236 6012
rect 8260 6010 8316 6012
rect 8340 6010 8396 6012
rect 8420 6010 8476 6012
rect 8180 5958 8226 6010
rect 8226 5958 8236 6010
rect 8260 5958 8290 6010
rect 8290 5958 8302 6010
rect 8302 5958 8316 6010
rect 8340 5958 8354 6010
rect 8354 5958 8366 6010
rect 8366 5958 8396 6010
rect 8420 5958 8430 6010
rect 8430 5958 8476 6010
rect 8180 5956 8236 5958
rect 8260 5956 8316 5958
rect 8340 5956 8396 5958
rect 8420 5956 8476 5958
rect 8180 4922 8236 4924
rect 8260 4922 8316 4924
rect 8340 4922 8396 4924
rect 8420 4922 8476 4924
rect 8180 4870 8226 4922
rect 8226 4870 8236 4922
rect 8260 4870 8290 4922
rect 8290 4870 8302 4922
rect 8302 4870 8316 4922
rect 8340 4870 8354 4922
rect 8354 4870 8366 4922
rect 8366 4870 8396 4922
rect 8420 4870 8430 4922
rect 8430 4870 8476 4922
rect 8180 4868 8236 4870
rect 8260 4868 8316 4870
rect 8340 4868 8396 4870
rect 8420 4868 8476 4870
rect 15404 26138 15460 26140
rect 15484 26138 15540 26140
rect 15564 26138 15620 26140
rect 15644 26138 15700 26140
rect 15404 26086 15450 26138
rect 15450 26086 15460 26138
rect 15484 26086 15514 26138
rect 15514 26086 15526 26138
rect 15526 26086 15540 26138
rect 15564 26086 15578 26138
rect 15578 26086 15590 26138
rect 15590 26086 15620 26138
rect 15644 26086 15654 26138
rect 15654 26086 15700 26138
rect 15404 26084 15460 26086
rect 15484 26084 15540 26086
rect 15564 26084 15620 26086
rect 15644 26084 15700 26086
rect 22628 33210 22684 33212
rect 22708 33210 22764 33212
rect 22788 33210 22844 33212
rect 22868 33210 22924 33212
rect 22628 33158 22674 33210
rect 22674 33158 22684 33210
rect 22708 33158 22738 33210
rect 22738 33158 22750 33210
rect 22750 33158 22764 33210
rect 22788 33158 22802 33210
rect 22802 33158 22814 33210
rect 22814 33158 22844 33210
rect 22868 33158 22878 33210
rect 22878 33158 22924 33210
rect 22628 33156 22684 33158
rect 22708 33156 22764 33158
rect 22788 33156 22844 33158
rect 22868 33156 22924 33158
rect 22628 32122 22684 32124
rect 22708 32122 22764 32124
rect 22788 32122 22844 32124
rect 22868 32122 22924 32124
rect 22628 32070 22674 32122
rect 22674 32070 22684 32122
rect 22708 32070 22738 32122
rect 22738 32070 22750 32122
rect 22750 32070 22764 32122
rect 22788 32070 22802 32122
rect 22802 32070 22814 32122
rect 22814 32070 22844 32122
rect 22868 32070 22878 32122
rect 22878 32070 22924 32122
rect 22628 32068 22684 32070
rect 22708 32068 22764 32070
rect 22788 32068 22844 32070
rect 22868 32068 22924 32070
rect 22628 31034 22684 31036
rect 22708 31034 22764 31036
rect 22788 31034 22844 31036
rect 22868 31034 22924 31036
rect 22628 30982 22674 31034
rect 22674 30982 22684 31034
rect 22708 30982 22738 31034
rect 22738 30982 22750 31034
rect 22750 30982 22764 31034
rect 22788 30982 22802 31034
rect 22802 30982 22814 31034
rect 22814 30982 22844 31034
rect 22868 30982 22878 31034
rect 22878 30982 22924 31034
rect 22628 30980 22684 30982
rect 22708 30980 22764 30982
rect 22788 30980 22844 30982
rect 22868 30980 22924 30982
rect 22628 29946 22684 29948
rect 22708 29946 22764 29948
rect 22788 29946 22844 29948
rect 22868 29946 22924 29948
rect 22628 29894 22674 29946
rect 22674 29894 22684 29946
rect 22708 29894 22738 29946
rect 22738 29894 22750 29946
rect 22750 29894 22764 29946
rect 22788 29894 22802 29946
rect 22802 29894 22814 29946
rect 22814 29894 22844 29946
rect 22868 29894 22878 29946
rect 22878 29894 22924 29946
rect 22628 29892 22684 29894
rect 22708 29892 22764 29894
rect 22788 29892 22844 29894
rect 22868 29892 22924 29894
rect 15404 25050 15460 25052
rect 15484 25050 15540 25052
rect 15564 25050 15620 25052
rect 15644 25050 15700 25052
rect 15404 24998 15450 25050
rect 15450 24998 15460 25050
rect 15484 24998 15514 25050
rect 15514 24998 15526 25050
rect 15526 24998 15540 25050
rect 15564 24998 15578 25050
rect 15578 24998 15590 25050
rect 15590 24998 15620 25050
rect 15644 24998 15654 25050
rect 15654 24998 15700 25050
rect 15404 24996 15460 24998
rect 15484 24996 15540 24998
rect 15564 24996 15620 24998
rect 15644 24996 15700 24998
rect 15404 23962 15460 23964
rect 15484 23962 15540 23964
rect 15564 23962 15620 23964
rect 15644 23962 15700 23964
rect 15404 23910 15450 23962
rect 15450 23910 15460 23962
rect 15484 23910 15514 23962
rect 15514 23910 15526 23962
rect 15526 23910 15540 23962
rect 15564 23910 15578 23962
rect 15578 23910 15590 23962
rect 15590 23910 15620 23962
rect 15644 23910 15654 23962
rect 15654 23910 15700 23962
rect 15404 23908 15460 23910
rect 15484 23908 15540 23910
rect 15564 23908 15620 23910
rect 15644 23908 15700 23910
rect 15404 22874 15460 22876
rect 15484 22874 15540 22876
rect 15564 22874 15620 22876
rect 15644 22874 15700 22876
rect 15404 22822 15450 22874
rect 15450 22822 15460 22874
rect 15484 22822 15514 22874
rect 15514 22822 15526 22874
rect 15526 22822 15540 22874
rect 15564 22822 15578 22874
rect 15578 22822 15590 22874
rect 15590 22822 15620 22874
rect 15644 22822 15654 22874
rect 15654 22822 15700 22874
rect 15404 22820 15460 22822
rect 15484 22820 15540 22822
rect 15564 22820 15620 22822
rect 15644 22820 15700 22822
rect 15404 21786 15460 21788
rect 15484 21786 15540 21788
rect 15564 21786 15620 21788
rect 15644 21786 15700 21788
rect 15404 21734 15450 21786
rect 15450 21734 15460 21786
rect 15484 21734 15514 21786
rect 15514 21734 15526 21786
rect 15526 21734 15540 21786
rect 15564 21734 15578 21786
rect 15578 21734 15590 21786
rect 15590 21734 15620 21786
rect 15644 21734 15654 21786
rect 15654 21734 15700 21786
rect 15404 21732 15460 21734
rect 15484 21732 15540 21734
rect 15564 21732 15620 21734
rect 15644 21732 15700 21734
rect 15404 20698 15460 20700
rect 15484 20698 15540 20700
rect 15564 20698 15620 20700
rect 15644 20698 15700 20700
rect 15404 20646 15450 20698
rect 15450 20646 15460 20698
rect 15484 20646 15514 20698
rect 15514 20646 15526 20698
rect 15526 20646 15540 20698
rect 15564 20646 15578 20698
rect 15578 20646 15590 20698
rect 15590 20646 15620 20698
rect 15644 20646 15654 20698
rect 15654 20646 15700 20698
rect 15404 20644 15460 20646
rect 15484 20644 15540 20646
rect 15564 20644 15620 20646
rect 15644 20644 15700 20646
rect 15842 20032 15898 20088
rect 14554 18128 14610 18184
rect 14094 16632 14150 16688
rect 15404 19610 15460 19612
rect 15484 19610 15540 19612
rect 15564 19610 15620 19612
rect 15644 19610 15700 19612
rect 15404 19558 15450 19610
rect 15450 19558 15460 19610
rect 15484 19558 15514 19610
rect 15514 19558 15526 19610
rect 15526 19558 15540 19610
rect 15564 19558 15578 19610
rect 15578 19558 15590 19610
rect 15590 19558 15620 19610
rect 15644 19558 15654 19610
rect 15654 19558 15700 19610
rect 15404 19556 15460 19558
rect 15484 19556 15540 19558
rect 15564 19556 15620 19558
rect 15644 19556 15700 19558
rect 14922 17176 14978 17232
rect 15404 18522 15460 18524
rect 15484 18522 15540 18524
rect 15564 18522 15620 18524
rect 15644 18522 15700 18524
rect 15404 18470 15450 18522
rect 15450 18470 15460 18522
rect 15484 18470 15514 18522
rect 15514 18470 15526 18522
rect 15526 18470 15540 18522
rect 15564 18470 15578 18522
rect 15578 18470 15590 18522
rect 15590 18470 15620 18522
rect 15644 18470 15654 18522
rect 15654 18470 15700 18522
rect 15404 18468 15460 18470
rect 15484 18468 15540 18470
rect 15564 18468 15620 18470
rect 15644 18468 15700 18470
rect 15106 17584 15162 17640
rect 17406 25236 17408 25256
rect 17408 25236 17460 25256
rect 17460 25236 17462 25256
rect 17406 25200 17462 25236
rect 17222 22616 17278 22672
rect 16578 19760 16634 19816
rect 16486 19624 16542 19680
rect 16026 18400 16082 18456
rect 15404 17434 15460 17436
rect 15484 17434 15540 17436
rect 15564 17434 15620 17436
rect 15644 17434 15700 17436
rect 15404 17382 15450 17434
rect 15450 17382 15460 17434
rect 15484 17382 15514 17434
rect 15514 17382 15526 17434
rect 15526 17382 15540 17434
rect 15564 17382 15578 17434
rect 15578 17382 15590 17434
rect 15590 17382 15620 17434
rect 15644 17382 15654 17434
rect 15654 17382 15700 17434
rect 15404 17380 15460 17382
rect 15484 17380 15540 17382
rect 15564 17380 15620 17382
rect 15644 17380 15700 17382
rect 15404 16346 15460 16348
rect 15484 16346 15540 16348
rect 15564 16346 15620 16348
rect 15644 16346 15700 16348
rect 15404 16294 15450 16346
rect 15450 16294 15460 16346
rect 15484 16294 15514 16346
rect 15514 16294 15526 16346
rect 15526 16294 15540 16346
rect 15564 16294 15578 16346
rect 15578 16294 15590 16346
rect 15590 16294 15620 16346
rect 15644 16294 15654 16346
rect 15654 16294 15700 16346
rect 15404 16292 15460 16294
rect 15484 16292 15540 16294
rect 15564 16292 15620 16294
rect 15644 16292 15700 16294
rect 15404 15258 15460 15260
rect 15484 15258 15540 15260
rect 15564 15258 15620 15260
rect 15644 15258 15700 15260
rect 15404 15206 15450 15258
rect 15450 15206 15460 15258
rect 15484 15206 15514 15258
rect 15514 15206 15526 15258
rect 15526 15206 15540 15258
rect 15564 15206 15578 15258
rect 15578 15206 15590 15258
rect 15590 15206 15620 15258
rect 15644 15206 15654 15258
rect 15654 15206 15700 15258
rect 15404 15204 15460 15206
rect 15484 15204 15540 15206
rect 15564 15204 15620 15206
rect 15644 15204 15700 15206
rect 15404 14170 15460 14172
rect 15484 14170 15540 14172
rect 15564 14170 15620 14172
rect 15644 14170 15700 14172
rect 15404 14118 15450 14170
rect 15450 14118 15460 14170
rect 15484 14118 15514 14170
rect 15514 14118 15526 14170
rect 15526 14118 15540 14170
rect 15564 14118 15578 14170
rect 15578 14118 15590 14170
rect 15590 14118 15620 14170
rect 15644 14118 15654 14170
rect 15654 14118 15700 14170
rect 15404 14116 15460 14118
rect 15484 14116 15540 14118
rect 15564 14116 15620 14118
rect 15644 14116 15700 14118
rect 15404 13082 15460 13084
rect 15484 13082 15540 13084
rect 15564 13082 15620 13084
rect 15644 13082 15700 13084
rect 15404 13030 15450 13082
rect 15450 13030 15460 13082
rect 15484 13030 15514 13082
rect 15514 13030 15526 13082
rect 15526 13030 15540 13082
rect 15564 13030 15578 13082
rect 15578 13030 15590 13082
rect 15590 13030 15620 13082
rect 15644 13030 15654 13082
rect 15654 13030 15700 13082
rect 15404 13028 15460 13030
rect 15484 13028 15540 13030
rect 15564 13028 15620 13030
rect 15644 13028 15700 13030
rect 15404 11994 15460 11996
rect 15484 11994 15540 11996
rect 15564 11994 15620 11996
rect 15644 11994 15700 11996
rect 15404 11942 15450 11994
rect 15450 11942 15460 11994
rect 15484 11942 15514 11994
rect 15514 11942 15526 11994
rect 15526 11942 15540 11994
rect 15564 11942 15578 11994
rect 15578 11942 15590 11994
rect 15590 11942 15620 11994
rect 15644 11942 15654 11994
rect 15654 11942 15700 11994
rect 15404 11940 15460 11942
rect 15484 11940 15540 11942
rect 15564 11940 15620 11942
rect 15644 11940 15700 11942
rect 16578 14320 16634 14376
rect 16394 12164 16450 12200
rect 16394 12144 16396 12164
rect 16396 12144 16448 12164
rect 16448 12144 16450 12164
rect 15404 10906 15460 10908
rect 15484 10906 15540 10908
rect 15564 10906 15620 10908
rect 15644 10906 15700 10908
rect 15404 10854 15450 10906
rect 15450 10854 15460 10906
rect 15484 10854 15514 10906
rect 15514 10854 15526 10906
rect 15526 10854 15540 10906
rect 15564 10854 15578 10906
rect 15578 10854 15590 10906
rect 15590 10854 15620 10906
rect 15644 10854 15654 10906
rect 15654 10854 15700 10906
rect 15404 10852 15460 10854
rect 15484 10852 15540 10854
rect 15564 10852 15620 10854
rect 15644 10852 15700 10854
rect 17222 16496 17278 16552
rect 17498 14900 17500 14920
rect 17500 14900 17552 14920
rect 17552 14900 17554 14920
rect 17498 14864 17554 14900
rect 17314 13232 17370 13288
rect 18050 23044 18106 23080
rect 18050 23024 18052 23044
rect 18052 23024 18104 23044
rect 18104 23024 18106 23044
rect 17774 17992 17830 18048
rect 18326 25200 18382 25256
rect 18418 23160 18474 23216
rect 18418 22500 18474 22536
rect 18418 22480 18420 22500
rect 18420 22480 18472 22500
rect 18472 22480 18474 22500
rect 18418 19896 18474 19952
rect 18142 13776 18198 13832
rect 8180 3834 8236 3836
rect 8260 3834 8316 3836
rect 8340 3834 8396 3836
rect 8420 3834 8476 3836
rect 8180 3782 8226 3834
rect 8226 3782 8236 3834
rect 8260 3782 8290 3834
rect 8290 3782 8302 3834
rect 8302 3782 8316 3834
rect 8340 3782 8354 3834
rect 8354 3782 8366 3834
rect 8366 3782 8396 3834
rect 8420 3782 8430 3834
rect 8430 3782 8476 3834
rect 8180 3780 8236 3782
rect 8260 3780 8316 3782
rect 8340 3780 8396 3782
rect 8420 3780 8476 3782
rect 8180 2746 8236 2748
rect 8260 2746 8316 2748
rect 8340 2746 8396 2748
rect 8420 2746 8476 2748
rect 8180 2694 8226 2746
rect 8226 2694 8236 2746
rect 8260 2694 8290 2746
rect 8290 2694 8302 2746
rect 8302 2694 8316 2746
rect 8340 2694 8354 2746
rect 8354 2694 8366 2746
rect 8366 2694 8396 2746
rect 8420 2694 8430 2746
rect 8430 2694 8476 2746
rect 8180 2692 8236 2694
rect 8260 2692 8316 2694
rect 8340 2692 8396 2694
rect 8420 2692 8476 2694
rect 15404 9818 15460 9820
rect 15484 9818 15540 9820
rect 15564 9818 15620 9820
rect 15644 9818 15700 9820
rect 15404 9766 15450 9818
rect 15450 9766 15460 9818
rect 15484 9766 15514 9818
rect 15514 9766 15526 9818
rect 15526 9766 15540 9818
rect 15564 9766 15578 9818
rect 15578 9766 15590 9818
rect 15590 9766 15620 9818
rect 15644 9766 15654 9818
rect 15654 9766 15700 9818
rect 15404 9764 15460 9766
rect 15484 9764 15540 9766
rect 15564 9764 15620 9766
rect 15644 9764 15700 9766
rect 18878 21800 18934 21856
rect 18694 18400 18750 18456
rect 18694 15988 18696 16008
rect 18696 15988 18748 16008
rect 18748 15988 18750 16008
rect 18694 15952 18750 15988
rect 19338 21972 19340 21992
rect 19340 21972 19392 21992
rect 19392 21972 19394 21992
rect 19338 21936 19394 21972
rect 19430 21664 19486 21720
rect 19246 18672 19302 18728
rect 19614 19796 19616 19816
rect 19616 19796 19668 19816
rect 19668 19796 19670 19816
rect 19614 19760 19670 19796
rect 19890 23704 19946 23760
rect 20534 24248 20590 24304
rect 20810 24656 20866 24712
rect 20718 23160 20774 23216
rect 21362 24148 21364 24168
rect 21364 24148 21416 24168
rect 21416 24148 21418 24168
rect 21362 24112 21418 24148
rect 21086 23568 21142 23624
rect 19890 19760 19946 19816
rect 18970 14456 19026 14512
rect 18326 12144 18382 12200
rect 21546 21020 21548 21040
rect 21548 21020 21600 21040
rect 21600 21020 21602 21040
rect 21546 20984 21602 21020
rect 19706 16224 19762 16280
rect 20074 15952 20130 16008
rect 19430 11600 19486 11656
rect 21178 17060 21234 17096
rect 21178 17040 21180 17060
rect 21180 17040 21232 17060
rect 21232 17040 21234 17060
rect 20902 15544 20958 15600
rect 20994 14048 21050 14104
rect 18418 9560 18474 9616
rect 15404 8730 15460 8732
rect 15484 8730 15540 8732
rect 15564 8730 15620 8732
rect 15644 8730 15700 8732
rect 15404 8678 15450 8730
rect 15450 8678 15460 8730
rect 15484 8678 15514 8730
rect 15514 8678 15526 8730
rect 15526 8678 15540 8730
rect 15564 8678 15578 8730
rect 15578 8678 15590 8730
rect 15590 8678 15620 8730
rect 15644 8678 15654 8730
rect 15654 8678 15700 8730
rect 15404 8676 15460 8678
rect 15484 8676 15540 8678
rect 15564 8676 15620 8678
rect 15644 8676 15700 8678
rect 15404 7642 15460 7644
rect 15484 7642 15540 7644
rect 15564 7642 15620 7644
rect 15644 7642 15700 7644
rect 15404 7590 15450 7642
rect 15450 7590 15460 7642
rect 15484 7590 15514 7642
rect 15514 7590 15526 7642
rect 15526 7590 15540 7642
rect 15564 7590 15578 7642
rect 15578 7590 15590 7642
rect 15590 7590 15620 7642
rect 15644 7590 15654 7642
rect 15654 7590 15700 7642
rect 15404 7588 15460 7590
rect 15484 7588 15540 7590
rect 15564 7588 15620 7590
rect 15644 7588 15700 7590
rect 15404 6554 15460 6556
rect 15484 6554 15540 6556
rect 15564 6554 15620 6556
rect 15644 6554 15700 6556
rect 15404 6502 15450 6554
rect 15450 6502 15460 6554
rect 15484 6502 15514 6554
rect 15514 6502 15526 6554
rect 15526 6502 15540 6554
rect 15564 6502 15578 6554
rect 15578 6502 15590 6554
rect 15590 6502 15620 6554
rect 15644 6502 15654 6554
rect 15654 6502 15700 6554
rect 15404 6500 15460 6502
rect 15484 6500 15540 6502
rect 15564 6500 15620 6502
rect 15644 6500 15700 6502
rect 15404 5466 15460 5468
rect 15484 5466 15540 5468
rect 15564 5466 15620 5468
rect 15644 5466 15700 5468
rect 15404 5414 15450 5466
rect 15450 5414 15460 5466
rect 15484 5414 15514 5466
rect 15514 5414 15526 5466
rect 15526 5414 15540 5466
rect 15564 5414 15578 5466
rect 15578 5414 15590 5466
rect 15590 5414 15620 5466
rect 15644 5414 15654 5466
rect 15654 5414 15700 5466
rect 15404 5412 15460 5414
rect 15484 5412 15540 5414
rect 15564 5412 15620 5414
rect 15644 5412 15700 5414
rect 15404 4378 15460 4380
rect 15484 4378 15540 4380
rect 15564 4378 15620 4380
rect 15644 4378 15700 4380
rect 15404 4326 15450 4378
rect 15450 4326 15460 4378
rect 15484 4326 15514 4378
rect 15514 4326 15526 4378
rect 15526 4326 15540 4378
rect 15564 4326 15578 4378
rect 15578 4326 15590 4378
rect 15590 4326 15620 4378
rect 15644 4326 15654 4378
rect 15654 4326 15700 4378
rect 15404 4324 15460 4326
rect 15484 4324 15540 4326
rect 15564 4324 15620 4326
rect 15644 4324 15700 4326
rect 15404 3290 15460 3292
rect 15484 3290 15540 3292
rect 15564 3290 15620 3292
rect 15644 3290 15700 3292
rect 15404 3238 15450 3290
rect 15450 3238 15460 3290
rect 15484 3238 15514 3290
rect 15514 3238 15526 3290
rect 15526 3238 15540 3290
rect 15564 3238 15578 3290
rect 15578 3238 15590 3290
rect 15590 3238 15620 3290
rect 15644 3238 15654 3290
rect 15654 3238 15700 3290
rect 15404 3236 15460 3238
rect 15484 3236 15540 3238
rect 15564 3236 15620 3238
rect 15644 3236 15700 3238
rect 21638 15000 21694 15056
rect 21178 8880 21234 8936
rect 22628 28858 22684 28860
rect 22708 28858 22764 28860
rect 22788 28858 22844 28860
rect 22868 28858 22924 28860
rect 22628 28806 22674 28858
rect 22674 28806 22684 28858
rect 22708 28806 22738 28858
rect 22738 28806 22750 28858
rect 22750 28806 22764 28858
rect 22788 28806 22802 28858
rect 22802 28806 22814 28858
rect 22814 28806 22844 28858
rect 22868 28806 22878 28858
rect 22878 28806 22924 28858
rect 22628 28804 22684 28806
rect 22708 28804 22764 28806
rect 22788 28804 22844 28806
rect 22868 28804 22924 28806
rect 22628 27770 22684 27772
rect 22708 27770 22764 27772
rect 22788 27770 22844 27772
rect 22868 27770 22924 27772
rect 22628 27718 22674 27770
rect 22674 27718 22684 27770
rect 22708 27718 22738 27770
rect 22738 27718 22750 27770
rect 22750 27718 22764 27770
rect 22788 27718 22802 27770
rect 22802 27718 22814 27770
rect 22814 27718 22844 27770
rect 22868 27718 22878 27770
rect 22878 27718 22924 27770
rect 22628 27716 22684 27718
rect 22708 27716 22764 27718
rect 22788 27716 22844 27718
rect 22868 27716 22924 27718
rect 22628 26682 22684 26684
rect 22708 26682 22764 26684
rect 22788 26682 22844 26684
rect 22868 26682 22924 26684
rect 22628 26630 22674 26682
rect 22674 26630 22684 26682
rect 22708 26630 22738 26682
rect 22738 26630 22750 26682
rect 22750 26630 22764 26682
rect 22788 26630 22802 26682
rect 22802 26630 22814 26682
rect 22814 26630 22844 26682
rect 22868 26630 22878 26682
rect 22878 26630 22924 26682
rect 22628 26628 22684 26630
rect 22708 26628 22764 26630
rect 22788 26628 22844 26630
rect 22868 26628 22924 26630
rect 22628 25594 22684 25596
rect 22708 25594 22764 25596
rect 22788 25594 22844 25596
rect 22868 25594 22924 25596
rect 22628 25542 22674 25594
rect 22674 25542 22684 25594
rect 22708 25542 22738 25594
rect 22738 25542 22750 25594
rect 22750 25542 22764 25594
rect 22788 25542 22802 25594
rect 22802 25542 22814 25594
rect 22814 25542 22844 25594
rect 22868 25542 22878 25594
rect 22878 25542 22924 25594
rect 22628 25540 22684 25542
rect 22708 25540 22764 25542
rect 22788 25540 22844 25542
rect 22868 25540 22924 25542
rect 22628 24506 22684 24508
rect 22708 24506 22764 24508
rect 22788 24506 22844 24508
rect 22868 24506 22924 24508
rect 22628 24454 22674 24506
rect 22674 24454 22684 24506
rect 22708 24454 22738 24506
rect 22738 24454 22750 24506
rect 22750 24454 22764 24506
rect 22788 24454 22802 24506
rect 22802 24454 22814 24506
rect 22814 24454 22844 24506
rect 22868 24454 22878 24506
rect 22878 24454 22924 24506
rect 22628 24452 22684 24454
rect 22708 24452 22764 24454
rect 22788 24452 22844 24454
rect 22868 24452 22924 24454
rect 22628 23418 22684 23420
rect 22708 23418 22764 23420
rect 22788 23418 22844 23420
rect 22868 23418 22924 23420
rect 22628 23366 22674 23418
rect 22674 23366 22684 23418
rect 22708 23366 22738 23418
rect 22738 23366 22750 23418
rect 22750 23366 22764 23418
rect 22788 23366 22802 23418
rect 22802 23366 22814 23418
rect 22814 23366 22844 23418
rect 22868 23366 22878 23418
rect 22878 23366 22924 23418
rect 22628 23364 22684 23366
rect 22708 23364 22764 23366
rect 22788 23364 22844 23366
rect 22868 23364 22924 23366
rect 22628 22330 22684 22332
rect 22708 22330 22764 22332
rect 22788 22330 22844 22332
rect 22868 22330 22924 22332
rect 22628 22278 22674 22330
rect 22674 22278 22684 22330
rect 22708 22278 22738 22330
rect 22738 22278 22750 22330
rect 22750 22278 22764 22330
rect 22788 22278 22802 22330
rect 22802 22278 22814 22330
rect 22814 22278 22844 22330
rect 22868 22278 22878 22330
rect 22878 22278 22924 22330
rect 22628 22276 22684 22278
rect 22708 22276 22764 22278
rect 22788 22276 22844 22278
rect 22868 22276 22924 22278
rect 22098 21936 22154 21992
rect 21822 21800 21878 21856
rect 22742 21972 22744 21992
rect 22744 21972 22796 21992
rect 22796 21972 22798 21992
rect 22742 21936 22798 21972
rect 22628 21242 22684 21244
rect 22708 21242 22764 21244
rect 22788 21242 22844 21244
rect 22868 21242 22924 21244
rect 22628 21190 22674 21242
rect 22674 21190 22684 21242
rect 22708 21190 22738 21242
rect 22738 21190 22750 21242
rect 22750 21190 22764 21242
rect 22788 21190 22802 21242
rect 22802 21190 22814 21242
rect 22814 21190 22844 21242
rect 22868 21190 22878 21242
rect 22878 21190 22924 21242
rect 22628 21188 22684 21190
rect 22708 21188 22764 21190
rect 22788 21188 22844 21190
rect 22868 21188 22924 21190
rect 22628 20154 22684 20156
rect 22708 20154 22764 20156
rect 22788 20154 22844 20156
rect 22868 20154 22924 20156
rect 22628 20102 22674 20154
rect 22674 20102 22684 20154
rect 22708 20102 22738 20154
rect 22738 20102 22750 20154
rect 22750 20102 22764 20154
rect 22788 20102 22802 20154
rect 22802 20102 22814 20154
rect 22814 20102 22844 20154
rect 22868 20102 22878 20154
rect 22878 20102 22924 20154
rect 22628 20100 22684 20102
rect 22708 20100 22764 20102
rect 22788 20100 22844 20102
rect 22868 20100 22924 20102
rect 22190 20032 22246 20088
rect 22190 18264 22246 18320
rect 21822 17312 21878 17368
rect 22006 14356 22008 14376
rect 22008 14356 22060 14376
rect 22060 14356 22062 14376
rect 22006 14320 22062 14356
rect 22628 19066 22684 19068
rect 22708 19066 22764 19068
rect 22788 19066 22844 19068
rect 22868 19066 22924 19068
rect 22628 19014 22674 19066
rect 22674 19014 22684 19066
rect 22708 19014 22738 19066
rect 22738 19014 22750 19066
rect 22750 19014 22764 19066
rect 22788 19014 22802 19066
rect 22802 19014 22814 19066
rect 22814 19014 22844 19066
rect 22868 19014 22878 19066
rect 22878 19014 22924 19066
rect 22628 19012 22684 19014
rect 22708 19012 22764 19014
rect 22788 19012 22844 19014
rect 22868 19012 22924 19014
rect 22374 18264 22430 18320
rect 22374 17992 22430 18048
rect 22628 17978 22684 17980
rect 22708 17978 22764 17980
rect 22788 17978 22844 17980
rect 22868 17978 22924 17980
rect 22628 17926 22674 17978
rect 22674 17926 22684 17978
rect 22708 17926 22738 17978
rect 22738 17926 22750 17978
rect 22750 17926 22764 17978
rect 22788 17926 22802 17978
rect 22802 17926 22814 17978
rect 22814 17926 22844 17978
rect 22868 17926 22878 17978
rect 22878 17926 22924 17978
rect 22628 17924 22684 17926
rect 22708 17924 22764 17926
rect 22788 17924 22844 17926
rect 22868 17924 22924 17926
rect 22628 16890 22684 16892
rect 22708 16890 22764 16892
rect 22788 16890 22844 16892
rect 22868 16890 22924 16892
rect 22628 16838 22674 16890
rect 22674 16838 22684 16890
rect 22708 16838 22738 16890
rect 22738 16838 22750 16890
rect 22750 16838 22764 16890
rect 22788 16838 22802 16890
rect 22802 16838 22814 16890
rect 22814 16838 22844 16890
rect 22868 16838 22878 16890
rect 22878 16838 22924 16890
rect 22628 16836 22684 16838
rect 22708 16836 22764 16838
rect 22788 16836 22844 16838
rect 22868 16836 22924 16838
rect 22628 15802 22684 15804
rect 22708 15802 22764 15804
rect 22788 15802 22844 15804
rect 22868 15802 22924 15804
rect 22628 15750 22674 15802
rect 22674 15750 22684 15802
rect 22708 15750 22738 15802
rect 22738 15750 22750 15802
rect 22750 15750 22764 15802
rect 22788 15750 22802 15802
rect 22802 15750 22814 15802
rect 22814 15750 22844 15802
rect 22868 15750 22878 15802
rect 22878 15750 22924 15802
rect 22628 15748 22684 15750
rect 22708 15748 22764 15750
rect 22788 15748 22844 15750
rect 22868 15748 22924 15750
rect 23938 22072 23994 22128
rect 37076 33210 37132 33212
rect 37156 33210 37212 33212
rect 37236 33210 37292 33212
rect 37316 33210 37372 33212
rect 37076 33158 37122 33210
rect 37122 33158 37132 33210
rect 37156 33158 37186 33210
rect 37186 33158 37198 33210
rect 37198 33158 37212 33210
rect 37236 33158 37250 33210
rect 37250 33158 37262 33210
rect 37262 33158 37292 33210
rect 37316 33158 37326 33210
rect 37326 33158 37372 33210
rect 37076 33156 37132 33158
rect 37156 33156 37212 33158
rect 37236 33156 37292 33158
rect 37316 33156 37372 33158
rect 29852 32666 29908 32668
rect 29932 32666 29988 32668
rect 30012 32666 30068 32668
rect 30092 32666 30148 32668
rect 29852 32614 29898 32666
rect 29898 32614 29908 32666
rect 29932 32614 29962 32666
rect 29962 32614 29974 32666
rect 29974 32614 29988 32666
rect 30012 32614 30026 32666
rect 30026 32614 30038 32666
rect 30038 32614 30068 32666
rect 30092 32614 30102 32666
rect 30102 32614 30148 32666
rect 29852 32612 29908 32614
rect 29932 32612 29988 32614
rect 30012 32612 30068 32614
rect 30092 32612 30148 32614
rect 29852 31578 29908 31580
rect 29932 31578 29988 31580
rect 30012 31578 30068 31580
rect 30092 31578 30148 31580
rect 29852 31526 29898 31578
rect 29898 31526 29908 31578
rect 29932 31526 29962 31578
rect 29962 31526 29974 31578
rect 29974 31526 29988 31578
rect 30012 31526 30026 31578
rect 30026 31526 30038 31578
rect 30038 31526 30068 31578
rect 30092 31526 30102 31578
rect 30102 31526 30148 31578
rect 29852 31524 29908 31526
rect 29932 31524 29988 31526
rect 30012 31524 30068 31526
rect 30092 31524 30148 31526
rect 29852 30490 29908 30492
rect 29932 30490 29988 30492
rect 30012 30490 30068 30492
rect 30092 30490 30148 30492
rect 29852 30438 29898 30490
rect 29898 30438 29908 30490
rect 29932 30438 29962 30490
rect 29962 30438 29974 30490
rect 29974 30438 29988 30490
rect 30012 30438 30026 30490
rect 30026 30438 30038 30490
rect 30038 30438 30068 30490
rect 30092 30438 30102 30490
rect 30102 30438 30148 30490
rect 29852 30436 29908 30438
rect 29932 30436 29988 30438
rect 30012 30436 30068 30438
rect 30092 30436 30148 30438
rect 29852 29402 29908 29404
rect 29932 29402 29988 29404
rect 30012 29402 30068 29404
rect 30092 29402 30148 29404
rect 29852 29350 29898 29402
rect 29898 29350 29908 29402
rect 29932 29350 29962 29402
rect 29962 29350 29974 29402
rect 29974 29350 29988 29402
rect 30012 29350 30026 29402
rect 30026 29350 30038 29402
rect 30038 29350 30068 29402
rect 30092 29350 30102 29402
rect 30102 29350 30148 29402
rect 29852 29348 29908 29350
rect 29932 29348 29988 29350
rect 30012 29348 30068 29350
rect 30092 29348 30148 29350
rect 26330 25356 26386 25392
rect 26330 25336 26332 25356
rect 26332 25336 26384 25356
rect 26384 25336 26386 25356
rect 24490 24812 24546 24848
rect 24490 24792 24492 24812
rect 24492 24792 24544 24812
rect 24544 24792 24546 24812
rect 24490 23044 24546 23080
rect 24490 23024 24492 23044
rect 24492 23024 24544 23044
rect 24544 23024 24546 23044
rect 24490 22072 24546 22128
rect 24490 21528 24546 21584
rect 24306 20576 24362 20632
rect 23294 17196 23350 17232
rect 23294 17176 23296 17196
rect 23296 17176 23348 17196
rect 23348 17176 23350 17196
rect 22628 14714 22684 14716
rect 22708 14714 22764 14716
rect 22788 14714 22844 14716
rect 22868 14714 22924 14716
rect 22628 14662 22674 14714
rect 22674 14662 22684 14714
rect 22708 14662 22738 14714
rect 22738 14662 22750 14714
rect 22750 14662 22764 14714
rect 22788 14662 22802 14714
rect 22802 14662 22814 14714
rect 22814 14662 22844 14714
rect 22868 14662 22878 14714
rect 22878 14662 22924 14714
rect 22628 14660 22684 14662
rect 22708 14660 22764 14662
rect 22788 14660 22844 14662
rect 22868 14660 22924 14662
rect 22628 13626 22684 13628
rect 22708 13626 22764 13628
rect 22788 13626 22844 13628
rect 22868 13626 22924 13628
rect 22628 13574 22674 13626
rect 22674 13574 22684 13626
rect 22708 13574 22738 13626
rect 22738 13574 22750 13626
rect 22750 13574 22764 13626
rect 22788 13574 22802 13626
rect 22802 13574 22814 13626
rect 22814 13574 22844 13626
rect 22868 13574 22878 13626
rect 22878 13574 22924 13626
rect 22628 13572 22684 13574
rect 22708 13572 22764 13574
rect 22788 13572 22844 13574
rect 22868 13572 22924 13574
rect 22628 12538 22684 12540
rect 22708 12538 22764 12540
rect 22788 12538 22844 12540
rect 22868 12538 22924 12540
rect 22628 12486 22674 12538
rect 22674 12486 22684 12538
rect 22708 12486 22738 12538
rect 22738 12486 22750 12538
rect 22750 12486 22764 12538
rect 22788 12486 22802 12538
rect 22802 12486 22814 12538
rect 22814 12486 22844 12538
rect 22868 12486 22878 12538
rect 22878 12486 22924 12538
rect 22628 12484 22684 12486
rect 22708 12484 22764 12486
rect 22788 12484 22844 12486
rect 22868 12484 22924 12486
rect 22282 12280 22338 12336
rect 23478 11756 23534 11792
rect 23478 11736 23480 11756
rect 23480 11736 23532 11756
rect 23532 11736 23534 11756
rect 21914 9968 21970 10024
rect 22628 11450 22684 11452
rect 22708 11450 22764 11452
rect 22788 11450 22844 11452
rect 22868 11450 22924 11452
rect 22628 11398 22674 11450
rect 22674 11398 22684 11450
rect 22708 11398 22738 11450
rect 22738 11398 22750 11450
rect 22750 11398 22764 11450
rect 22788 11398 22802 11450
rect 22802 11398 22814 11450
rect 22814 11398 22844 11450
rect 22868 11398 22878 11450
rect 22878 11398 22924 11450
rect 22628 11396 22684 11398
rect 22708 11396 22764 11398
rect 22788 11396 22844 11398
rect 22868 11396 22924 11398
rect 25226 23024 25282 23080
rect 25042 21664 25098 21720
rect 25502 23160 25558 23216
rect 26146 21664 26202 21720
rect 27434 24112 27490 24168
rect 26882 23060 26884 23080
rect 26884 23060 26936 23080
rect 26936 23060 26938 23080
rect 26882 23024 26938 23060
rect 27066 21528 27122 21584
rect 28262 20576 28318 20632
rect 27250 19624 27306 19680
rect 22628 10362 22684 10364
rect 22708 10362 22764 10364
rect 22788 10362 22844 10364
rect 22868 10362 22924 10364
rect 22628 10310 22674 10362
rect 22674 10310 22684 10362
rect 22708 10310 22738 10362
rect 22738 10310 22750 10362
rect 22750 10310 22764 10362
rect 22788 10310 22802 10362
rect 22802 10310 22814 10362
rect 22814 10310 22844 10362
rect 22868 10310 22878 10362
rect 22878 10310 22924 10362
rect 22628 10308 22684 10310
rect 22708 10308 22764 10310
rect 22788 10308 22844 10310
rect 22868 10308 22924 10310
rect 26146 12180 26148 12200
rect 26148 12180 26200 12200
rect 26200 12180 26202 12200
rect 26146 12144 26202 12180
rect 27342 18264 27398 18320
rect 26790 17040 26846 17096
rect 26882 12280 26938 12336
rect 27618 14048 27674 14104
rect 22628 9274 22684 9276
rect 22708 9274 22764 9276
rect 22788 9274 22844 9276
rect 22868 9274 22924 9276
rect 22628 9222 22674 9274
rect 22674 9222 22684 9274
rect 22708 9222 22738 9274
rect 22738 9222 22750 9274
rect 22750 9222 22764 9274
rect 22788 9222 22802 9274
rect 22802 9222 22814 9274
rect 22814 9222 22844 9274
rect 22868 9222 22878 9274
rect 22878 9222 22924 9274
rect 22628 9220 22684 9222
rect 22708 9220 22764 9222
rect 22788 9220 22844 9222
rect 22868 9220 22924 9222
rect 22628 8186 22684 8188
rect 22708 8186 22764 8188
rect 22788 8186 22844 8188
rect 22868 8186 22924 8188
rect 22628 8134 22674 8186
rect 22674 8134 22684 8186
rect 22708 8134 22738 8186
rect 22738 8134 22750 8186
rect 22750 8134 22764 8186
rect 22788 8134 22802 8186
rect 22802 8134 22814 8186
rect 22814 8134 22844 8186
rect 22868 8134 22878 8186
rect 22878 8134 22924 8186
rect 22628 8132 22684 8134
rect 22708 8132 22764 8134
rect 22788 8132 22844 8134
rect 22868 8132 22924 8134
rect 27802 7812 27858 7848
rect 27802 7792 27804 7812
rect 27804 7792 27856 7812
rect 27856 7792 27858 7812
rect 22628 7098 22684 7100
rect 22708 7098 22764 7100
rect 22788 7098 22844 7100
rect 22868 7098 22924 7100
rect 22628 7046 22674 7098
rect 22674 7046 22684 7098
rect 22708 7046 22738 7098
rect 22738 7046 22750 7098
rect 22750 7046 22764 7098
rect 22788 7046 22802 7098
rect 22802 7046 22814 7098
rect 22814 7046 22844 7098
rect 22868 7046 22878 7098
rect 22878 7046 22924 7098
rect 22628 7044 22684 7046
rect 22708 7044 22764 7046
rect 22788 7044 22844 7046
rect 22868 7044 22924 7046
rect 22628 6010 22684 6012
rect 22708 6010 22764 6012
rect 22788 6010 22844 6012
rect 22868 6010 22924 6012
rect 22628 5958 22674 6010
rect 22674 5958 22684 6010
rect 22708 5958 22738 6010
rect 22738 5958 22750 6010
rect 22750 5958 22764 6010
rect 22788 5958 22802 6010
rect 22802 5958 22814 6010
rect 22814 5958 22844 6010
rect 22868 5958 22878 6010
rect 22878 5958 22924 6010
rect 22628 5956 22684 5958
rect 22708 5956 22764 5958
rect 22788 5956 22844 5958
rect 22868 5956 22924 5958
rect 22628 4922 22684 4924
rect 22708 4922 22764 4924
rect 22788 4922 22844 4924
rect 22868 4922 22924 4924
rect 22628 4870 22674 4922
rect 22674 4870 22684 4922
rect 22708 4870 22738 4922
rect 22738 4870 22750 4922
rect 22750 4870 22764 4922
rect 22788 4870 22802 4922
rect 22802 4870 22814 4922
rect 22814 4870 22844 4922
rect 22868 4870 22878 4922
rect 22878 4870 22924 4922
rect 22628 4868 22684 4870
rect 22708 4868 22764 4870
rect 22788 4868 22844 4870
rect 22868 4868 22924 4870
rect 24858 4564 24860 4584
rect 24860 4564 24912 4584
rect 24912 4564 24914 4584
rect 24858 4528 24914 4564
rect 22628 3834 22684 3836
rect 22708 3834 22764 3836
rect 22788 3834 22844 3836
rect 22868 3834 22924 3836
rect 22628 3782 22674 3834
rect 22674 3782 22684 3834
rect 22708 3782 22738 3834
rect 22738 3782 22750 3834
rect 22750 3782 22764 3834
rect 22788 3782 22802 3834
rect 22802 3782 22814 3834
rect 22814 3782 22844 3834
rect 22868 3782 22878 3834
rect 22878 3782 22924 3834
rect 22628 3780 22684 3782
rect 22708 3780 22764 3782
rect 22788 3780 22844 3782
rect 22868 3780 22924 3782
rect 28354 17312 28410 17368
rect 28814 15000 28870 15056
rect 28262 7404 28318 7440
rect 28262 7384 28264 7404
rect 28264 7384 28316 7404
rect 28316 7384 28318 7404
rect 28814 6976 28870 7032
rect 29852 28314 29908 28316
rect 29932 28314 29988 28316
rect 30012 28314 30068 28316
rect 30092 28314 30148 28316
rect 29852 28262 29898 28314
rect 29898 28262 29908 28314
rect 29932 28262 29962 28314
rect 29962 28262 29974 28314
rect 29974 28262 29988 28314
rect 30012 28262 30026 28314
rect 30026 28262 30038 28314
rect 30038 28262 30068 28314
rect 30092 28262 30102 28314
rect 30102 28262 30148 28314
rect 29852 28260 29908 28262
rect 29932 28260 29988 28262
rect 30012 28260 30068 28262
rect 30092 28260 30148 28262
rect 29852 27226 29908 27228
rect 29932 27226 29988 27228
rect 30012 27226 30068 27228
rect 30092 27226 30148 27228
rect 29852 27174 29898 27226
rect 29898 27174 29908 27226
rect 29932 27174 29962 27226
rect 29962 27174 29974 27226
rect 29974 27174 29988 27226
rect 30012 27174 30026 27226
rect 30026 27174 30038 27226
rect 30038 27174 30068 27226
rect 30092 27174 30102 27226
rect 30102 27174 30148 27226
rect 29852 27172 29908 27174
rect 29932 27172 29988 27174
rect 30012 27172 30068 27174
rect 30092 27172 30148 27174
rect 29852 26138 29908 26140
rect 29932 26138 29988 26140
rect 30012 26138 30068 26140
rect 30092 26138 30148 26140
rect 29852 26086 29898 26138
rect 29898 26086 29908 26138
rect 29932 26086 29962 26138
rect 29962 26086 29974 26138
rect 29974 26086 29988 26138
rect 30012 26086 30026 26138
rect 30026 26086 30038 26138
rect 30038 26086 30068 26138
rect 30092 26086 30102 26138
rect 30102 26086 30148 26138
rect 29852 26084 29908 26086
rect 29932 26084 29988 26086
rect 30012 26084 30068 26086
rect 30092 26084 30148 26086
rect 29852 25050 29908 25052
rect 29932 25050 29988 25052
rect 30012 25050 30068 25052
rect 30092 25050 30148 25052
rect 29852 24998 29898 25050
rect 29898 24998 29908 25050
rect 29932 24998 29962 25050
rect 29962 24998 29974 25050
rect 29974 24998 29988 25050
rect 30012 24998 30026 25050
rect 30026 24998 30038 25050
rect 30038 24998 30068 25050
rect 30092 24998 30102 25050
rect 30102 24998 30148 25050
rect 29852 24996 29908 24998
rect 29932 24996 29988 24998
rect 30012 24996 30068 24998
rect 30092 24996 30148 24998
rect 29852 23962 29908 23964
rect 29932 23962 29988 23964
rect 30012 23962 30068 23964
rect 30092 23962 30148 23964
rect 29852 23910 29898 23962
rect 29898 23910 29908 23962
rect 29932 23910 29962 23962
rect 29962 23910 29974 23962
rect 29974 23910 29988 23962
rect 30012 23910 30026 23962
rect 30026 23910 30038 23962
rect 30038 23910 30068 23962
rect 30092 23910 30102 23962
rect 30102 23910 30148 23962
rect 29852 23908 29908 23910
rect 29932 23908 29988 23910
rect 30012 23908 30068 23910
rect 30092 23908 30148 23910
rect 29852 22874 29908 22876
rect 29932 22874 29988 22876
rect 30012 22874 30068 22876
rect 30092 22874 30148 22876
rect 29852 22822 29898 22874
rect 29898 22822 29908 22874
rect 29932 22822 29962 22874
rect 29962 22822 29974 22874
rect 29974 22822 29988 22874
rect 30012 22822 30026 22874
rect 30026 22822 30038 22874
rect 30038 22822 30068 22874
rect 30092 22822 30102 22874
rect 30102 22822 30148 22874
rect 29852 22820 29908 22822
rect 29932 22820 29988 22822
rect 30012 22820 30068 22822
rect 30092 22820 30148 22822
rect 29366 21412 29422 21448
rect 29366 21392 29368 21412
rect 29368 21392 29420 21412
rect 29420 21392 29422 21412
rect 29852 21786 29908 21788
rect 29932 21786 29988 21788
rect 30012 21786 30068 21788
rect 30092 21786 30148 21788
rect 29852 21734 29898 21786
rect 29898 21734 29908 21786
rect 29932 21734 29962 21786
rect 29962 21734 29974 21786
rect 29974 21734 29988 21786
rect 30012 21734 30026 21786
rect 30026 21734 30038 21786
rect 30038 21734 30068 21786
rect 30092 21734 30102 21786
rect 30102 21734 30148 21786
rect 29852 21732 29908 21734
rect 29932 21732 29988 21734
rect 30012 21732 30068 21734
rect 30092 21732 30148 21734
rect 29852 20698 29908 20700
rect 29932 20698 29988 20700
rect 30012 20698 30068 20700
rect 30092 20698 30148 20700
rect 29852 20646 29898 20698
rect 29898 20646 29908 20698
rect 29932 20646 29962 20698
rect 29962 20646 29974 20698
rect 29974 20646 29988 20698
rect 30012 20646 30026 20698
rect 30026 20646 30038 20698
rect 30038 20646 30068 20698
rect 30092 20646 30102 20698
rect 30102 20646 30148 20698
rect 29852 20644 29908 20646
rect 29932 20644 29988 20646
rect 30012 20644 30068 20646
rect 30092 20644 30148 20646
rect 29852 19610 29908 19612
rect 29932 19610 29988 19612
rect 30012 19610 30068 19612
rect 30092 19610 30148 19612
rect 29852 19558 29898 19610
rect 29898 19558 29908 19610
rect 29932 19558 29962 19610
rect 29962 19558 29974 19610
rect 29974 19558 29988 19610
rect 30012 19558 30026 19610
rect 30026 19558 30038 19610
rect 30038 19558 30068 19610
rect 30092 19558 30102 19610
rect 30102 19558 30148 19610
rect 29852 19556 29908 19558
rect 29932 19556 29988 19558
rect 30012 19556 30068 19558
rect 30092 19556 30148 19558
rect 29852 18522 29908 18524
rect 29932 18522 29988 18524
rect 30012 18522 30068 18524
rect 30092 18522 30148 18524
rect 29852 18470 29898 18522
rect 29898 18470 29908 18522
rect 29932 18470 29962 18522
rect 29962 18470 29974 18522
rect 29974 18470 29988 18522
rect 30012 18470 30026 18522
rect 30026 18470 30038 18522
rect 30038 18470 30068 18522
rect 30092 18470 30102 18522
rect 30102 18470 30148 18522
rect 29852 18468 29908 18470
rect 29932 18468 29988 18470
rect 30012 18468 30068 18470
rect 30092 18468 30148 18470
rect 28998 15408 29054 15464
rect 29550 16224 29606 16280
rect 29852 17434 29908 17436
rect 29932 17434 29988 17436
rect 30012 17434 30068 17436
rect 30092 17434 30148 17436
rect 29852 17382 29898 17434
rect 29898 17382 29908 17434
rect 29932 17382 29962 17434
rect 29962 17382 29974 17434
rect 29974 17382 29988 17434
rect 30012 17382 30026 17434
rect 30026 17382 30038 17434
rect 30038 17382 30068 17434
rect 30092 17382 30102 17434
rect 30102 17382 30148 17434
rect 29852 17380 29908 17382
rect 29932 17380 29988 17382
rect 30012 17380 30068 17382
rect 30092 17380 30148 17382
rect 29852 16346 29908 16348
rect 29932 16346 29988 16348
rect 30012 16346 30068 16348
rect 30092 16346 30148 16348
rect 29852 16294 29898 16346
rect 29898 16294 29908 16346
rect 29932 16294 29962 16346
rect 29962 16294 29974 16346
rect 29974 16294 29988 16346
rect 30012 16294 30026 16346
rect 30026 16294 30038 16346
rect 30038 16294 30068 16346
rect 30092 16294 30102 16346
rect 30102 16294 30148 16346
rect 29852 16292 29908 16294
rect 29932 16292 29988 16294
rect 30012 16292 30068 16294
rect 30092 16292 30148 16294
rect 29642 15952 29698 16008
rect 29852 15258 29908 15260
rect 29932 15258 29988 15260
rect 30012 15258 30068 15260
rect 30092 15258 30148 15260
rect 29852 15206 29898 15258
rect 29898 15206 29908 15258
rect 29932 15206 29962 15258
rect 29962 15206 29974 15258
rect 29974 15206 29988 15258
rect 30012 15206 30026 15258
rect 30026 15206 30038 15258
rect 30038 15206 30068 15258
rect 30092 15206 30102 15258
rect 30102 15206 30148 15258
rect 29852 15204 29908 15206
rect 29932 15204 29988 15206
rect 30012 15204 30068 15206
rect 30092 15204 30148 15206
rect 29852 14170 29908 14172
rect 29932 14170 29988 14172
rect 30012 14170 30068 14172
rect 30092 14170 30148 14172
rect 29852 14118 29898 14170
rect 29898 14118 29908 14170
rect 29932 14118 29962 14170
rect 29962 14118 29974 14170
rect 29974 14118 29988 14170
rect 30012 14118 30026 14170
rect 30026 14118 30038 14170
rect 30038 14118 30068 14170
rect 30092 14118 30102 14170
rect 30102 14118 30148 14170
rect 29852 14116 29908 14118
rect 29932 14116 29988 14118
rect 30012 14116 30068 14118
rect 30092 14116 30148 14118
rect 31206 17604 31262 17640
rect 31206 17584 31208 17604
rect 31208 17584 31260 17604
rect 31260 17584 31262 17604
rect 30930 13912 30986 13968
rect 29852 13082 29908 13084
rect 29932 13082 29988 13084
rect 30012 13082 30068 13084
rect 30092 13082 30148 13084
rect 29852 13030 29898 13082
rect 29898 13030 29908 13082
rect 29932 13030 29962 13082
rect 29962 13030 29974 13082
rect 29974 13030 29988 13082
rect 30012 13030 30026 13082
rect 30026 13030 30038 13082
rect 30038 13030 30068 13082
rect 30092 13030 30102 13082
rect 30102 13030 30148 13082
rect 29852 13028 29908 13030
rect 29932 13028 29988 13030
rect 30012 13028 30068 13030
rect 30092 13028 30148 13030
rect 29826 12860 29828 12880
rect 29828 12860 29880 12880
rect 29880 12860 29882 12880
rect 29826 12824 29882 12860
rect 29852 11994 29908 11996
rect 29932 11994 29988 11996
rect 30012 11994 30068 11996
rect 30092 11994 30148 11996
rect 29852 11942 29898 11994
rect 29898 11942 29908 11994
rect 29932 11942 29962 11994
rect 29962 11942 29974 11994
rect 29974 11942 29988 11994
rect 30012 11942 30026 11994
rect 30026 11942 30038 11994
rect 30038 11942 30068 11994
rect 30092 11942 30102 11994
rect 30102 11942 30148 11994
rect 29852 11940 29908 11942
rect 29932 11940 29988 11942
rect 30012 11940 30068 11942
rect 30092 11940 30148 11942
rect 29852 10906 29908 10908
rect 29932 10906 29988 10908
rect 30012 10906 30068 10908
rect 30092 10906 30148 10908
rect 29852 10854 29898 10906
rect 29898 10854 29908 10906
rect 29932 10854 29962 10906
rect 29962 10854 29974 10906
rect 29974 10854 29988 10906
rect 30012 10854 30026 10906
rect 30026 10854 30038 10906
rect 30038 10854 30068 10906
rect 30092 10854 30102 10906
rect 30102 10854 30148 10906
rect 29852 10852 29908 10854
rect 29932 10852 29988 10854
rect 30012 10852 30068 10854
rect 30092 10852 30148 10854
rect 30378 11600 30434 11656
rect 30286 9832 30342 9888
rect 29852 9818 29908 9820
rect 29932 9818 29988 9820
rect 30012 9818 30068 9820
rect 30092 9818 30148 9820
rect 29852 9766 29898 9818
rect 29898 9766 29908 9818
rect 29932 9766 29962 9818
rect 29962 9766 29974 9818
rect 29974 9766 29988 9818
rect 30012 9766 30026 9818
rect 30026 9766 30038 9818
rect 30038 9766 30068 9818
rect 30092 9766 30102 9818
rect 30102 9766 30148 9818
rect 29852 9764 29908 9766
rect 29932 9764 29988 9766
rect 30012 9764 30068 9766
rect 30092 9764 30148 9766
rect 29734 9016 29790 9072
rect 29852 8730 29908 8732
rect 29932 8730 29988 8732
rect 30012 8730 30068 8732
rect 30092 8730 30148 8732
rect 29852 8678 29898 8730
rect 29898 8678 29908 8730
rect 29932 8678 29962 8730
rect 29962 8678 29974 8730
rect 29974 8678 29988 8730
rect 30012 8678 30026 8730
rect 30026 8678 30038 8730
rect 30038 8678 30068 8730
rect 30092 8678 30102 8730
rect 30102 8678 30148 8730
rect 29852 8676 29908 8678
rect 29932 8676 29988 8678
rect 30012 8676 30068 8678
rect 30092 8676 30148 8678
rect 29852 7642 29908 7644
rect 29932 7642 29988 7644
rect 30012 7642 30068 7644
rect 30092 7642 30148 7644
rect 29852 7590 29898 7642
rect 29898 7590 29908 7642
rect 29932 7590 29962 7642
rect 29962 7590 29974 7642
rect 29974 7590 29988 7642
rect 30012 7590 30026 7642
rect 30026 7590 30038 7642
rect 30038 7590 30068 7642
rect 30092 7590 30102 7642
rect 30102 7590 30148 7642
rect 29852 7588 29908 7590
rect 29932 7588 29988 7590
rect 30012 7588 30068 7590
rect 30092 7588 30148 7590
rect 30470 10104 30526 10160
rect 30930 11620 30986 11656
rect 30930 11600 30932 11620
rect 30932 11600 30984 11620
rect 30984 11600 30986 11620
rect 32034 17584 32090 17640
rect 37076 32122 37132 32124
rect 37156 32122 37212 32124
rect 37236 32122 37292 32124
rect 37316 32122 37372 32124
rect 37076 32070 37122 32122
rect 37122 32070 37132 32122
rect 37156 32070 37186 32122
rect 37186 32070 37198 32122
rect 37198 32070 37212 32122
rect 37236 32070 37250 32122
rect 37250 32070 37262 32122
rect 37262 32070 37292 32122
rect 37316 32070 37326 32122
rect 37326 32070 37372 32122
rect 37076 32068 37132 32070
rect 37156 32068 37212 32070
rect 37236 32068 37292 32070
rect 37316 32068 37372 32070
rect 37076 31034 37132 31036
rect 37156 31034 37212 31036
rect 37236 31034 37292 31036
rect 37316 31034 37372 31036
rect 37076 30982 37122 31034
rect 37122 30982 37132 31034
rect 37156 30982 37186 31034
rect 37186 30982 37198 31034
rect 37198 30982 37212 31034
rect 37236 30982 37250 31034
rect 37250 30982 37262 31034
rect 37262 30982 37292 31034
rect 37316 30982 37326 31034
rect 37326 30982 37372 31034
rect 37076 30980 37132 30982
rect 37156 30980 37212 30982
rect 37236 30980 37292 30982
rect 37316 30980 37372 30982
rect 37076 29946 37132 29948
rect 37156 29946 37212 29948
rect 37236 29946 37292 29948
rect 37316 29946 37372 29948
rect 37076 29894 37122 29946
rect 37122 29894 37132 29946
rect 37156 29894 37186 29946
rect 37186 29894 37198 29946
rect 37198 29894 37212 29946
rect 37236 29894 37250 29946
rect 37250 29894 37262 29946
rect 37262 29894 37292 29946
rect 37316 29894 37326 29946
rect 37326 29894 37372 29946
rect 37076 29892 37132 29894
rect 37156 29892 37212 29894
rect 37236 29892 37292 29894
rect 37316 29892 37372 29894
rect 37076 28858 37132 28860
rect 37156 28858 37212 28860
rect 37236 28858 37292 28860
rect 37316 28858 37372 28860
rect 37076 28806 37122 28858
rect 37122 28806 37132 28858
rect 37156 28806 37186 28858
rect 37186 28806 37198 28858
rect 37198 28806 37212 28858
rect 37236 28806 37250 28858
rect 37250 28806 37262 28858
rect 37262 28806 37292 28858
rect 37316 28806 37326 28858
rect 37326 28806 37372 28858
rect 37076 28804 37132 28806
rect 37156 28804 37212 28806
rect 37236 28804 37292 28806
rect 37316 28804 37372 28806
rect 33598 23704 33654 23760
rect 32954 22480 33010 22536
rect 33598 18692 33654 18728
rect 33598 18672 33600 18692
rect 33600 18672 33652 18692
rect 33652 18672 33654 18692
rect 32126 16088 32182 16144
rect 37076 27770 37132 27772
rect 37156 27770 37212 27772
rect 37236 27770 37292 27772
rect 37316 27770 37372 27772
rect 37076 27718 37122 27770
rect 37122 27718 37132 27770
rect 37156 27718 37186 27770
rect 37186 27718 37198 27770
rect 37198 27718 37212 27770
rect 37236 27718 37250 27770
rect 37250 27718 37262 27770
rect 37262 27718 37292 27770
rect 37316 27718 37326 27770
rect 37326 27718 37372 27770
rect 37076 27716 37132 27718
rect 37156 27716 37212 27718
rect 37236 27716 37292 27718
rect 37316 27716 37372 27718
rect 34058 16632 34114 16688
rect 29852 6554 29908 6556
rect 29932 6554 29988 6556
rect 30012 6554 30068 6556
rect 30092 6554 30148 6556
rect 29852 6502 29898 6554
rect 29898 6502 29908 6554
rect 29932 6502 29962 6554
rect 29962 6502 29974 6554
rect 29974 6502 29988 6554
rect 30012 6502 30026 6554
rect 30026 6502 30038 6554
rect 30038 6502 30068 6554
rect 30092 6502 30102 6554
rect 30102 6502 30148 6554
rect 29852 6500 29908 6502
rect 29932 6500 29988 6502
rect 30012 6500 30068 6502
rect 30092 6500 30148 6502
rect 29852 5466 29908 5468
rect 29932 5466 29988 5468
rect 30012 5466 30068 5468
rect 30092 5466 30148 5468
rect 29852 5414 29898 5466
rect 29898 5414 29908 5466
rect 29932 5414 29962 5466
rect 29962 5414 29974 5466
rect 29974 5414 29988 5466
rect 30012 5414 30026 5466
rect 30026 5414 30038 5466
rect 30038 5414 30068 5466
rect 30092 5414 30102 5466
rect 30102 5414 30148 5466
rect 29852 5412 29908 5414
rect 29932 5412 29988 5414
rect 30012 5412 30068 5414
rect 30092 5412 30148 5414
rect 31666 9832 31722 9888
rect 30930 8492 30986 8528
rect 30930 8472 30932 8492
rect 30932 8472 30984 8492
rect 30984 8472 30986 8492
rect 31114 8064 31170 8120
rect 30562 6976 30618 7032
rect 31114 6976 31170 7032
rect 29852 4378 29908 4380
rect 29932 4378 29988 4380
rect 30012 4378 30068 4380
rect 30092 4378 30148 4380
rect 29852 4326 29898 4378
rect 29898 4326 29908 4378
rect 29932 4326 29962 4378
rect 29962 4326 29974 4378
rect 29974 4326 29988 4378
rect 30012 4326 30026 4378
rect 30026 4326 30038 4378
rect 30038 4326 30068 4378
rect 30092 4326 30102 4378
rect 30102 4326 30148 4378
rect 29852 4324 29908 4326
rect 29932 4324 29988 4326
rect 30012 4324 30068 4326
rect 30092 4324 30148 4326
rect 32770 9016 32826 9072
rect 31758 8064 31814 8120
rect 31666 7964 31668 7984
rect 31668 7964 31720 7984
rect 31720 7964 31722 7984
rect 31666 7928 31722 7964
rect 31574 6976 31630 7032
rect 31574 6860 31630 6896
rect 31574 6840 31576 6860
rect 31576 6840 31628 6860
rect 31628 6840 31630 6860
rect 37076 26682 37132 26684
rect 37156 26682 37212 26684
rect 37236 26682 37292 26684
rect 37316 26682 37372 26684
rect 37076 26630 37122 26682
rect 37122 26630 37132 26682
rect 37156 26630 37186 26682
rect 37186 26630 37198 26682
rect 37198 26630 37212 26682
rect 37236 26630 37250 26682
rect 37250 26630 37262 26682
rect 37262 26630 37292 26682
rect 37316 26630 37326 26682
rect 37326 26630 37372 26682
rect 37076 26628 37132 26630
rect 37156 26628 37212 26630
rect 37236 26628 37292 26630
rect 37316 26628 37372 26630
rect 37076 25594 37132 25596
rect 37156 25594 37212 25596
rect 37236 25594 37292 25596
rect 37316 25594 37372 25596
rect 37076 25542 37122 25594
rect 37122 25542 37132 25594
rect 37156 25542 37186 25594
rect 37186 25542 37198 25594
rect 37198 25542 37212 25594
rect 37236 25542 37250 25594
rect 37250 25542 37262 25594
rect 37262 25542 37292 25594
rect 37316 25542 37326 25594
rect 37326 25542 37372 25594
rect 37076 25540 37132 25542
rect 37156 25540 37212 25542
rect 37236 25540 37292 25542
rect 37316 25540 37372 25542
rect 37370 24692 37372 24712
rect 37372 24692 37424 24712
rect 37424 24692 37426 24712
rect 37370 24656 37426 24692
rect 37076 24506 37132 24508
rect 37156 24506 37212 24508
rect 37236 24506 37292 24508
rect 37316 24506 37372 24508
rect 37076 24454 37122 24506
rect 37122 24454 37132 24506
rect 37156 24454 37186 24506
rect 37186 24454 37198 24506
rect 37198 24454 37212 24506
rect 37236 24454 37250 24506
rect 37250 24454 37262 24506
rect 37262 24454 37292 24506
rect 37316 24454 37326 24506
rect 37326 24454 37372 24506
rect 37076 24452 37132 24454
rect 37156 24452 37212 24454
rect 37236 24452 37292 24454
rect 37316 24452 37372 24454
rect 37076 23418 37132 23420
rect 37156 23418 37212 23420
rect 37236 23418 37292 23420
rect 37316 23418 37372 23420
rect 37076 23366 37122 23418
rect 37122 23366 37132 23418
rect 37156 23366 37186 23418
rect 37186 23366 37198 23418
rect 37198 23366 37212 23418
rect 37236 23366 37250 23418
rect 37250 23366 37262 23418
rect 37262 23366 37292 23418
rect 37316 23366 37326 23418
rect 37326 23366 37372 23418
rect 37076 23364 37132 23366
rect 37156 23364 37212 23366
rect 37236 23364 37292 23366
rect 37316 23364 37372 23366
rect 37076 22330 37132 22332
rect 37156 22330 37212 22332
rect 37236 22330 37292 22332
rect 37316 22330 37372 22332
rect 37076 22278 37122 22330
rect 37122 22278 37132 22330
rect 37156 22278 37186 22330
rect 37186 22278 37198 22330
rect 37198 22278 37212 22330
rect 37236 22278 37250 22330
rect 37250 22278 37262 22330
rect 37262 22278 37292 22330
rect 37316 22278 37326 22330
rect 37326 22278 37372 22330
rect 37076 22276 37132 22278
rect 37156 22276 37212 22278
rect 37236 22276 37292 22278
rect 37316 22276 37372 22278
rect 36726 20984 36782 21040
rect 37076 21242 37132 21244
rect 37156 21242 37212 21244
rect 37236 21242 37292 21244
rect 37316 21242 37372 21244
rect 37076 21190 37122 21242
rect 37122 21190 37132 21242
rect 37156 21190 37186 21242
rect 37186 21190 37198 21242
rect 37198 21190 37212 21242
rect 37236 21190 37250 21242
rect 37250 21190 37262 21242
rect 37262 21190 37292 21242
rect 37316 21190 37326 21242
rect 37326 21190 37372 21242
rect 37076 21188 37132 21190
rect 37156 21188 37212 21190
rect 37236 21188 37292 21190
rect 37316 21188 37372 21190
rect 37076 20154 37132 20156
rect 37156 20154 37212 20156
rect 37236 20154 37292 20156
rect 37316 20154 37372 20156
rect 37076 20102 37122 20154
rect 37122 20102 37132 20154
rect 37156 20102 37186 20154
rect 37186 20102 37198 20154
rect 37198 20102 37212 20154
rect 37236 20102 37250 20154
rect 37250 20102 37262 20154
rect 37262 20102 37292 20154
rect 37316 20102 37326 20154
rect 37326 20102 37372 20154
rect 37076 20100 37132 20102
rect 37156 20100 37212 20102
rect 37236 20100 37292 20102
rect 37316 20100 37372 20102
rect 37076 19066 37132 19068
rect 37156 19066 37212 19068
rect 37236 19066 37292 19068
rect 37316 19066 37372 19068
rect 37076 19014 37122 19066
rect 37122 19014 37132 19066
rect 37156 19014 37186 19066
rect 37186 19014 37198 19066
rect 37198 19014 37212 19066
rect 37236 19014 37250 19066
rect 37250 19014 37262 19066
rect 37262 19014 37292 19066
rect 37316 19014 37326 19066
rect 37326 19014 37372 19066
rect 37076 19012 37132 19014
rect 37156 19012 37212 19014
rect 37236 19012 37292 19014
rect 37316 19012 37372 19014
rect 37076 17978 37132 17980
rect 37156 17978 37212 17980
rect 37236 17978 37292 17980
rect 37316 17978 37372 17980
rect 37076 17926 37122 17978
rect 37122 17926 37132 17978
rect 37156 17926 37186 17978
rect 37186 17926 37198 17978
rect 37198 17926 37212 17978
rect 37236 17926 37250 17978
rect 37250 17926 37262 17978
rect 37262 17926 37292 17978
rect 37316 17926 37326 17978
rect 37326 17926 37372 17978
rect 37076 17924 37132 17926
rect 37156 17924 37212 17926
rect 37236 17924 37292 17926
rect 37316 17924 37372 17926
rect 37076 16890 37132 16892
rect 37156 16890 37212 16892
rect 37236 16890 37292 16892
rect 37316 16890 37372 16892
rect 37076 16838 37122 16890
rect 37122 16838 37132 16890
rect 37156 16838 37186 16890
rect 37186 16838 37198 16890
rect 37198 16838 37212 16890
rect 37236 16838 37250 16890
rect 37250 16838 37262 16890
rect 37262 16838 37292 16890
rect 37316 16838 37326 16890
rect 37326 16838 37372 16890
rect 37076 16836 37132 16838
rect 37156 16836 37212 16838
rect 37236 16836 37292 16838
rect 37316 16836 37372 16838
rect 37076 15802 37132 15804
rect 37156 15802 37212 15804
rect 37236 15802 37292 15804
rect 37316 15802 37372 15804
rect 37076 15750 37122 15802
rect 37122 15750 37132 15802
rect 37156 15750 37186 15802
rect 37186 15750 37198 15802
rect 37198 15750 37212 15802
rect 37236 15750 37250 15802
rect 37250 15750 37262 15802
rect 37262 15750 37292 15802
rect 37316 15750 37326 15802
rect 37326 15750 37372 15802
rect 37076 15748 37132 15750
rect 37156 15748 37212 15750
rect 37236 15748 37292 15750
rect 37316 15748 37372 15750
rect 37076 14714 37132 14716
rect 37156 14714 37212 14716
rect 37236 14714 37292 14716
rect 37316 14714 37372 14716
rect 37076 14662 37122 14714
rect 37122 14662 37132 14714
rect 37156 14662 37186 14714
rect 37186 14662 37198 14714
rect 37198 14662 37212 14714
rect 37236 14662 37250 14714
rect 37250 14662 37262 14714
rect 37262 14662 37292 14714
rect 37316 14662 37326 14714
rect 37326 14662 37372 14714
rect 37076 14660 37132 14662
rect 37156 14660 37212 14662
rect 37236 14660 37292 14662
rect 37316 14660 37372 14662
rect 37076 13626 37132 13628
rect 37156 13626 37212 13628
rect 37236 13626 37292 13628
rect 37316 13626 37372 13628
rect 37076 13574 37122 13626
rect 37122 13574 37132 13626
rect 37156 13574 37186 13626
rect 37186 13574 37198 13626
rect 37198 13574 37212 13626
rect 37236 13574 37250 13626
rect 37250 13574 37262 13626
rect 37262 13574 37292 13626
rect 37316 13574 37326 13626
rect 37326 13574 37372 13626
rect 37076 13572 37132 13574
rect 37156 13572 37212 13574
rect 37236 13572 37292 13574
rect 37316 13572 37372 13574
rect 37076 12538 37132 12540
rect 37156 12538 37212 12540
rect 37236 12538 37292 12540
rect 37316 12538 37372 12540
rect 37076 12486 37122 12538
rect 37122 12486 37132 12538
rect 37156 12486 37186 12538
rect 37186 12486 37198 12538
rect 37198 12486 37212 12538
rect 37236 12486 37250 12538
rect 37250 12486 37262 12538
rect 37262 12486 37292 12538
rect 37316 12486 37326 12538
rect 37326 12486 37372 12538
rect 37076 12484 37132 12486
rect 37156 12484 37212 12486
rect 37236 12484 37292 12486
rect 37316 12484 37372 12486
rect 33046 7404 33102 7440
rect 33046 7384 33048 7404
rect 33048 7384 33100 7404
rect 33100 7384 33102 7404
rect 29852 3290 29908 3292
rect 29932 3290 29988 3292
rect 30012 3290 30068 3292
rect 30092 3290 30148 3292
rect 29852 3238 29898 3290
rect 29898 3238 29908 3290
rect 29932 3238 29962 3290
rect 29962 3238 29974 3290
rect 29974 3238 29988 3290
rect 30012 3238 30026 3290
rect 30026 3238 30038 3290
rect 30038 3238 30068 3290
rect 30092 3238 30102 3290
rect 30102 3238 30148 3290
rect 29852 3236 29908 3238
rect 29932 3236 29988 3238
rect 30012 3236 30068 3238
rect 30092 3236 30148 3238
rect 33690 7828 33692 7848
rect 33692 7828 33744 7848
rect 33744 7828 33746 7848
rect 33690 7792 33746 7828
rect 37076 11450 37132 11452
rect 37156 11450 37212 11452
rect 37236 11450 37292 11452
rect 37316 11450 37372 11452
rect 37076 11398 37122 11450
rect 37122 11398 37132 11450
rect 37156 11398 37186 11450
rect 37186 11398 37198 11450
rect 37198 11398 37212 11450
rect 37236 11398 37250 11450
rect 37250 11398 37262 11450
rect 37262 11398 37292 11450
rect 37316 11398 37326 11450
rect 37326 11398 37372 11450
rect 37076 11396 37132 11398
rect 37156 11396 37212 11398
rect 37236 11396 37292 11398
rect 37316 11396 37372 11398
rect 38014 21392 38070 21448
rect 39210 19780 39266 19816
rect 39210 19760 39212 19780
rect 39212 19760 39264 19780
rect 39264 19760 39266 19780
rect 38842 18128 38898 18184
rect 38106 17620 38108 17640
rect 38108 17620 38160 17640
rect 38160 17620 38162 17640
rect 38106 17584 38162 17620
rect 38658 17176 38714 17232
rect 38566 15680 38622 15736
rect 37738 10668 37794 10704
rect 37738 10648 37740 10668
rect 37740 10648 37792 10668
rect 37792 10648 37794 10668
rect 37076 10362 37132 10364
rect 37156 10362 37212 10364
rect 37236 10362 37292 10364
rect 37316 10362 37372 10364
rect 37076 10310 37122 10362
rect 37122 10310 37132 10362
rect 37156 10310 37186 10362
rect 37186 10310 37198 10362
rect 37198 10310 37212 10362
rect 37236 10310 37250 10362
rect 37250 10310 37262 10362
rect 37262 10310 37292 10362
rect 37316 10310 37326 10362
rect 37326 10310 37372 10362
rect 37076 10308 37132 10310
rect 37156 10308 37212 10310
rect 37236 10308 37292 10310
rect 37316 10308 37372 10310
rect 36910 10124 36966 10160
rect 36910 10104 36912 10124
rect 36912 10104 36964 10124
rect 36964 10104 36966 10124
rect 37076 9274 37132 9276
rect 37156 9274 37212 9276
rect 37236 9274 37292 9276
rect 37316 9274 37372 9276
rect 37076 9222 37122 9274
rect 37122 9222 37132 9274
rect 37156 9222 37186 9274
rect 37186 9222 37198 9274
rect 37198 9222 37212 9274
rect 37236 9222 37250 9274
rect 37250 9222 37262 9274
rect 37262 9222 37292 9274
rect 37316 9222 37326 9274
rect 37326 9222 37372 9274
rect 37076 9220 37132 9222
rect 37156 9220 37212 9222
rect 37236 9220 37292 9222
rect 37316 9220 37372 9222
rect 37076 8186 37132 8188
rect 37156 8186 37212 8188
rect 37236 8186 37292 8188
rect 37316 8186 37372 8188
rect 37076 8134 37122 8186
rect 37122 8134 37132 8186
rect 37156 8134 37186 8186
rect 37186 8134 37198 8186
rect 37198 8134 37212 8186
rect 37236 8134 37250 8186
rect 37250 8134 37262 8186
rect 37262 8134 37292 8186
rect 37316 8134 37326 8186
rect 37326 8134 37372 8186
rect 37076 8132 37132 8134
rect 37156 8132 37212 8134
rect 37236 8132 37292 8134
rect 37316 8132 37372 8134
rect 37076 7098 37132 7100
rect 37156 7098 37212 7100
rect 37236 7098 37292 7100
rect 37316 7098 37372 7100
rect 37076 7046 37122 7098
rect 37122 7046 37132 7098
rect 37156 7046 37186 7098
rect 37186 7046 37198 7098
rect 37198 7046 37212 7098
rect 37236 7046 37250 7098
rect 37250 7046 37262 7098
rect 37262 7046 37292 7098
rect 37316 7046 37326 7098
rect 37326 7046 37372 7098
rect 37076 7044 37132 7046
rect 37156 7044 37212 7046
rect 37236 7044 37292 7046
rect 37316 7044 37372 7046
rect 37076 6010 37132 6012
rect 37156 6010 37212 6012
rect 37236 6010 37292 6012
rect 37316 6010 37372 6012
rect 37076 5958 37122 6010
rect 37122 5958 37132 6010
rect 37156 5958 37186 6010
rect 37186 5958 37198 6010
rect 37198 5958 37212 6010
rect 37236 5958 37250 6010
rect 37250 5958 37262 6010
rect 37262 5958 37292 6010
rect 37316 5958 37326 6010
rect 37326 5958 37372 6010
rect 37076 5956 37132 5958
rect 37156 5956 37212 5958
rect 37236 5956 37292 5958
rect 37316 5956 37372 5958
rect 37076 4922 37132 4924
rect 37156 4922 37212 4924
rect 37236 4922 37292 4924
rect 37316 4922 37372 4924
rect 37076 4870 37122 4922
rect 37122 4870 37132 4922
rect 37156 4870 37186 4922
rect 37186 4870 37198 4922
rect 37198 4870 37212 4922
rect 37236 4870 37250 4922
rect 37250 4870 37262 4922
rect 37262 4870 37292 4922
rect 37316 4870 37326 4922
rect 37326 4870 37372 4922
rect 37076 4868 37132 4870
rect 37156 4868 37212 4870
rect 37236 4868 37292 4870
rect 37316 4868 37372 4870
rect 37076 3834 37132 3836
rect 37156 3834 37212 3836
rect 37236 3834 37292 3836
rect 37316 3834 37372 3836
rect 37076 3782 37122 3834
rect 37122 3782 37132 3834
rect 37156 3782 37186 3834
rect 37186 3782 37198 3834
rect 37198 3782 37212 3834
rect 37236 3782 37250 3834
rect 37250 3782 37262 3834
rect 37262 3782 37292 3834
rect 37316 3782 37326 3834
rect 37326 3782 37372 3834
rect 37076 3780 37132 3782
rect 37156 3780 37212 3782
rect 37236 3780 37292 3782
rect 37316 3780 37372 3782
rect 22628 2746 22684 2748
rect 22708 2746 22764 2748
rect 22788 2746 22844 2748
rect 22868 2746 22924 2748
rect 22628 2694 22674 2746
rect 22674 2694 22684 2746
rect 22708 2694 22738 2746
rect 22738 2694 22750 2746
rect 22750 2694 22764 2746
rect 22788 2694 22802 2746
rect 22802 2694 22814 2746
rect 22814 2694 22844 2746
rect 22868 2694 22878 2746
rect 22878 2694 22924 2746
rect 22628 2692 22684 2694
rect 22708 2692 22764 2694
rect 22788 2692 22844 2694
rect 22868 2692 22924 2694
rect 37076 2746 37132 2748
rect 37156 2746 37212 2748
rect 37236 2746 37292 2748
rect 37316 2746 37372 2748
rect 37076 2694 37122 2746
rect 37122 2694 37132 2746
rect 37156 2694 37186 2746
rect 37186 2694 37198 2746
rect 37198 2694 37212 2746
rect 37236 2694 37250 2746
rect 37250 2694 37262 2746
rect 37262 2694 37292 2746
rect 37316 2694 37326 2746
rect 37326 2694 37372 2746
rect 37076 2692 37132 2694
rect 37156 2692 37212 2694
rect 37236 2692 37292 2694
rect 37316 2692 37372 2694
rect 38106 11092 38108 11112
rect 38108 11092 38160 11112
rect 38160 11092 38162 11112
rect 38106 11056 38162 11092
rect 39118 15680 39174 15736
rect 41786 19916 41842 19952
rect 41786 19896 41788 19916
rect 41788 19896 41840 19916
rect 41840 19896 41842 19916
rect 43350 18128 43406 18184
rect 41602 15680 41658 15736
rect 38474 10648 38530 10704
rect 38658 9968 38714 10024
rect 38658 8608 38714 8664
rect 38290 6840 38346 6896
rect 39026 7928 39082 7984
rect 39762 8472 39818 8528
rect 39854 8336 39910 8392
rect 39670 8200 39726 8256
rect 40866 8608 40922 8664
rect 51524 33210 51580 33212
rect 51604 33210 51660 33212
rect 51684 33210 51740 33212
rect 51764 33210 51820 33212
rect 51524 33158 51570 33210
rect 51570 33158 51580 33210
rect 51604 33158 51634 33210
rect 51634 33158 51646 33210
rect 51646 33158 51660 33210
rect 51684 33158 51698 33210
rect 51698 33158 51710 33210
rect 51710 33158 51740 33210
rect 51764 33158 51774 33210
rect 51774 33158 51820 33210
rect 51524 33156 51580 33158
rect 51604 33156 51660 33158
rect 51684 33156 51740 33158
rect 51764 33156 51820 33158
rect 44300 32666 44356 32668
rect 44380 32666 44436 32668
rect 44460 32666 44516 32668
rect 44540 32666 44596 32668
rect 44300 32614 44346 32666
rect 44346 32614 44356 32666
rect 44380 32614 44410 32666
rect 44410 32614 44422 32666
rect 44422 32614 44436 32666
rect 44460 32614 44474 32666
rect 44474 32614 44486 32666
rect 44486 32614 44516 32666
rect 44540 32614 44550 32666
rect 44550 32614 44596 32666
rect 44300 32612 44356 32614
rect 44380 32612 44436 32614
rect 44460 32612 44516 32614
rect 44540 32612 44596 32614
rect 51524 32122 51580 32124
rect 51604 32122 51660 32124
rect 51684 32122 51740 32124
rect 51764 32122 51820 32124
rect 51524 32070 51570 32122
rect 51570 32070 51580 32122
rect 51604 32070 51634 32122
rect 51634 32070 51646 32122
rect 51646 32070 51660 32122
rect 51684 32070 51698 32122
rect 51698 32070 51710 32122
rect 51710 32070 51740 32122
rect 51764 32070 51774 32122
rect 51774 32070 51820 32122
rect 51524 32068 51580 32070
rect 51604 32068 51660 32070
rect 51684 32068 51740 32070
rect 51764 32068 51820 32070
rect 44300 31578 44356 31580
rect 44380 31578 44436 31580
rect 44460 31578 44516 31580
rect 44540 31578 44596 31580
rect 44300 31526 44346 31578
rect 44346 31526 44356 31578
rect 44380 31526 44410 31578
rect 44410 31526 44422 31578
rect 44422 31526 44436 31578
rect 44460 31526 44474 31578
rect 44474 31526 44486 31578
rect 44486 31526 44516 31578
rect 44540 31526 44550 31578
rect 44550 31526 44596 31578
rect 44300 31524 44356 31526
rect 44380 31524 44436 31526
rect 44460 31524 44516 31526
rect 44540 31524 44596 31526
rect 44300 30490 44356 30492
rect 44380 30490 44436 30492
rect 44460 30490 44516 30492
rect 44540 30490 44596 30492
rect 44300 30438 44346 30490
rect 44346 30438 44356 30490
rect 44380 30438 44410 30490
rect 44410 30438 44422 30490
rect 44422 30438 44436 30490
rect 44460 30438 44474 30490
rect 44474 30438 44486 30490
rect 44486 30438 44516 30490
rect 44540 30438 44550 30490
rect 44550 30438 44596 30490
rect 44300 30436 44356 30438
rect 44380 30436 44436 30438
rect 44460 30436 44516 30438
rect 44540 30436 44596 30438
rect 44300 29402 44356 29404
rect 44380 29402 44436 29404
rect 44460 29402 44516 29404
rect 44540 29402 44596 29404
rect 44300 29350 44346 29402
rect 44346 29350 44356 29402
rect 44380 29350 44410 29402
rect 44410 29350 44422 29402
rect 44422 29350 44436 29402
rect 44460 29350 44474 29402
rect 44474 29350 44486 29402
rect 44486 29350 44516 29402
rect 44540 29350 44550 29402
rect 44550 29350 44596 29402
rect 44300 29348 44356 29350
rect 44380 29348 44436 29350
rect 44460 29348 44516 29350
rect 44540 29348 44596 29350
rect 44300 28314 44356 28316
rect 44380 28314 44436 28316
rect 44460 28314 44516 28316
rect 44540 28314 44596 28316
rect 44300 28262 44346 28314
rect 44346 28262 44356 28314
rect 44380 28262 44410 28314
rect 44410 28262 44422 28314
rect 44422 28262 44436 28314
rect 44460 28262 44474 28314
rect 44474 28262 44486 28314
rect 44486 28262 44516 28314
rect 44540 28262 44550 28314
rect 44550 28262 44596 28314
rect 44300 28260 44356 28262
rect 44380 28260 44436 28262
rect 44460 28260 44516 28262
rect 44540 28260 44596 28262
rect 51524 31034 51580 31036
rect 51604 31034 51660 31036
rect 51684 31034 51740 31036
rect 51764 31034 51820 31036
rect 51524 30982 51570 31034
rect 51570 30982 51580 31034
rect 51604 30982 51634 31034
rect 51634 30982 51646 31034
rect 51646 30982 51660 31034
rect 51684 30982 51698 31034
rect 51698 30982 51710 31034
rect 51710 30982 51740 31034
rect 51764 30982 51774 31034
rect 51774 30982 51820 31034
rect 51524 30980 51580 30982
rect 51604 30980 51660 30982
rect 51684 30980 51740 30982
rect 51764 30980 51820 30982
rect 51524 29946 51580 29948
rect 51604 29946 51660 29948
rect 51684 29946 51740 29948
rect 51764 29946 51820 29948
rect 51524 29894 51570 29946
rect 51570 29894 51580 29946
rect 51604 29894 51634 29946
rect 51634 29894 51646 29946
rect 51646 29894 51660 29946
rect 51684 29894 51698 29946
rect 51698 29894 51710 29946
rect 51710 29894 51740 29946
rect 51764 29894 51774 29946
rect 51774 29894 51820 29946
rect 51524 29892 51580 29894
rect 51604 29892 51660 29894
rect 51684 29892 51740 29894
rect 51764 29892 51820 29894
rect 51524 28858 51580 28860
rect 51604 28858 51660 28860
rect 51684 28858 51740 28860
rect 51764 28858 51820 28860
rect 51524 28806 51570 28858
rect 51570 28806 51580 28858
rect 51604 28806 51634 28858
rect 51634 28806 51646 28858
rect 51646 28806 51660 28858
rect 51684 28806 51698 28858
rect 51698 28806 51710 28858
rect 51710 28806 51740 28858
rect 51764 28806 51774 28858
rect 51774 28806 51820 28858
rect 51524 28804 51580 28806
rect 51604 28804 51660 28806
rect 51684 28804 51740 28806
rect 51764 28804 51820 28806
rect 51524 27770 51580 27772
rect 51604 27770 51660 27772
rect 51684 27770 51740 27772
rect 51764 27770 51820 27772
rect 51524 27718 51570 27770
rect 51570 27718 51580 27770
rect 51604 27718 51634 27770
rect 51634 27718 51646 27770
rect 51646 27718 51660 27770
rect 51684 27718 51698 27770
rect 51698 27718 51710 27770
rect 51710 27718 51740 27770
rect 51764 27718 51774 27770
rect 51774 27718 51820 27770
rect 51524 27716 51580 27718
rect 51604 27716 51660 27718
rect 51684 27716 51740 27718
rect 51764 27716 51820 27718
rect 44300 27226 44356 27228
rect 44380 27226 44436 27228
rect 44460 27226 44516 27228
rect 44540 27226 44596 27228
rect 44300 27174 44346 27226
rect 44346 27174 44356 27226
rect 44380 27174 44410 27226
rect 44410 27174 44422 27226
rect 44422 27174 44436 27226
rect 44460 27174 44474 27226
rect 44474 27174 44486 27226
rect 44486 27174 44516 27226
rect 44540 27174 44550 27226
rect 44550 27174 44596 27226
rect 44300 27172 44356 27174
rect 44380 27172 44436 27174
rect 44460 27172 44516 27174
rect 44540 27172 44596 27174
rect 51524 26682 51580 26684
rect 51604 26682 51660 26684
rect 51684 26682 51740 26684
rect 51764 26682 51820 26684
rect 51524 26630 51570 26682
rect 51570 26630 51580 26682
rect 51604 26630 51634 26682
rect 51634 26630 51646 26682
rect 51646 26630 51660 26682
rect 51684 26630 51698 26682
rect 51698 26630 51710 26682
rect 51710 26630 51740 26682
rect 51764 26630 51774 26682
rect 51774 26630 51820 26682
rect 51524 26628 51580 26630
rect 51604 26628 51660 26630
rect 51684 26628 51740 26630
rect 51764 26628 51820 26630
rect 44300 26138 44356 26140
rect 44380 26138 44436 26140
rect 44460 26138 44516 26140
rect 44540 26138 44596 26140
rect 44300 26086 44346 26138
rect 44346 26086 44356 26138
rect 44380 26086 44410 26138
rect 44410 26086 44422 26138
rect 44422 26086 44436 26138
rect 44460 26086 44474 26138
rect 44474 26086 44486 26138
rect 44486 26086 44516 26138
rect 44540 26086 44550 26138
rect 44550 26086 44596 26138
rect 44300 26084 44356 26086
rect 44380 26084 44436 26086
rect 44460 26084 44516 26086
rect 44540 26084 44596 26086
rect 51524 25594 51580 25596
rect 51604 25594 51660 25596
rect 51684 25594 51740 25596
rect 51764 25594 51820 25596
rect 51524 25542 51570 25594
rect 51570 25542 51580 25594
rect 51604 25542 51634 25594
rect 51634 25542 51646 25594
rect 51646 25542 51660 25594
rect 51684 25542 51698 25594
rect 51698 25542 51710 25594
rect 51710 25542 51740 25594
rect 51764 25542 51774 25594
rect 51774 25542 51820 25594
rect 51524 25540 51580 25542
rect 51604 25540 51660 25542
rect 51684 25540 51740 25542
rect 51764 25540 51820 25542
rect 44300 25050 44356 25052
rect 44380 25050 44436 25052
rect 44460 25050 44516 25052
rect 44540 25050 44596 25052
rect 44300 24998 44346 25050
rect 44346 24998 44356 25050
rect 44380 24998 44410 25050
rect 44410 24998 44422 25050
rect 44422 24998 44436 25050
rect 44460 24998 44474 25050
rect 44474 24998 44486 25050
rect 44486 24998 44516 25050
rect 44540 24998 44550 25050
rect 44550 24998 44596 25050
rect 44300 24996 44356 24998
rect 44380 24996 44436 24998
rect 44460 24996 44516 24998
rect 44540 24996 44596 24998
rect 51524 24506 51580 24508
rect 51604 24506 51660 24508
rect 51684 24506 51740 24508
rect 51764 24506 51820 24508
rect 51524 24454 51570 24506
rect 51570 24454 51580 24506
rect 51604 24454 51634 24506
rect 51634 24454 51646 24506
rect 51646 24454 51660 24506
rect 51684 24454 51698 24506
rect 51698 24454 51710 24506
rect 51710 24454 51740 24506
rect 51764 24454 51774 24506
rect 51774 24454 51820 24506
rect 51524 24452 51580 24454
rect 51604 24452 51660 24454
rect 51684 24452 51740 24454
rect 51764 24452 51820 24454
rect 44300 23962 44356 23964
rect 44380 23962 44436 23964
rect 44460 23962 44516 23964
rect 44540 23962 44596 23964
rect 44300 23910 44346 23962
rect 44346 23910 44356 23962
rect 44380 23910 44410 23962
rect 44410 23910 44422 23962
rect 44422 23910 44436 23962
rect 44460 23910 44474 23962
rect 44474 23910 44486 23962
rect 44486 23910 44516 23962
rect 44540 23910 44550 23962
rect 44550 23910 44596 23962
rect 44300 23908 44356 23910
rect 44380 23908 44436 23910
rect 44460 23908 44516 23910
rect 44540 23908 44596 23910
rect 44300 22874 44356 22876
rect 44380 22874 44436 22876
rect 44460 22874 44516 22876
rect 44540 22874 44596 22876
rect 44300 22822 44346 22874
rect 44346 22822 44356 22874
rect 44380 22822 44410 22874
rect 44410 22822 44422 22874
rect 44422 22822 44436 22874
rect 44460 22822 44474 22874
rect 44474 22822 44486 22874
rect 44486 22822 44516 22874
rect 44540 22822 44550 22874
rect 44550 22822 44596 22874
rect 44300 22820 44356 22822
rect 44380 22820 44436 22822
rect 44460 22820 44516 22822
rect 44540 22820 44596 22822
rect 44300 21786 44356 21788
rect 44380 21786 44436 21788
rect 44460 21786 44516 21788
rect 44540 21786 44596 21788
rect 44300 21734 44346 21786
rect 44346 21734 44356 21786
rect 44380 21734 44410 21786
rect 44410 21734 44422 21786
rect 44422 21734 44436 21786
rect 44460 21734 44474 21786
rect 44474 21734 44486 21786
rect 44486 21734 44516 21786
rect 44540 21734 44550 21786
rect 44550 21734 44596 21786
rect 44300 21732 44356 21734
rect 44380 21732 44436 21734
rect 44460 21732 44516 21734
rect 44540 21732 44596 21734
rect 44300 20698 44356 20700
rect 44380 20698 44436 20700
rect 44460 20698 44516 20700
rect 44540 20698 44596 20700
rect 44300 20646 44346 20698
rect 44346 20646 44356 20698
rect 44380 20646 44410 20698
rect 44410 20646 44422 20698
rect 44422 20646 44436 20698
rect 44460 20646 44474 20698
rect 44474 20646 44486 20698
rect 44486 20646 44516 20698
rect 44540 20646 44550 20698
rect 44550 20646 44596 20698
rect 44300 20644 44356 20646
rect 44380 20644 44436 20646
rect 44460 20644 44516 20646
rect 44540 20644 44596 20646
rect 44300 19610 44356 19612
rect 44380 19610 44436 19612
rect 44460 19610 44516 19612
rect 44540 19610 44596 19612
rect 44300 19558 44346 19610
rect 44346 19558 44356 19610
rect 44380 19558 44410 19610
rect 44410 19558 44422 19610
rect 44422 19558 44436 19610
rect 44460 19558 44474 19610
rect 44474 19558 44486 19610
rect 44486 19558 44516 19610
rect 44540 19558 44550 19610
rect 44550 19558 44596 19610
rect 44300 19556 44356 19558
rect 44380 19556 44436 19558
rect 44460 19556 44516 19558
rect 44540 19556 44596 19558
rect 44300 18522 44356 18524
rect 44380 18522 44436 18524
rect 44460 18522 44516 18524
rect 44540 18522 44596 18524
rect 44300 18470 44346 18522
rect 44346 18470 44356 18522
rect 44380 18470 44410 18522
rect 44410 18470 44422 18522
rect 44422 18470 44436 18522
rect 44460 18470 44474 18522
rect 44474 18470 44486 18522
rect 44486 18470 44516 18522
rect 44540 18470 44550 18522
rect 44550 18470 44596 18522
rect 44300 18468 44356 18470
rect 44380 18468 44436 18470
rect 44460 18468 44516 18470
rect 44540 18468 44596 18470
rect 44300 17434 44356 17436
rect 44380 17434 44436 17436
rect 44460 17434 44516 17436
rect 44540 17434 44596 17436
rect 44300 17382 44346 17434
rect 44346 17382 44356 17434
rect 44380 17382 44410 17434
rect 44410 17382 44422 17434
rect 44422 17382 44436 17434
rect 44460 17382 44474 17434
rect 44474 17382 44486 17434
rect 44486 17382 44516 17434
rect 44540 17382 44550 17434
rect 44550 17382 44596 17434
rect 44300 17380 44356 17382
rect 44380 17380 44436 17382
rect 44460 17380 44516 17382
rect 44540 17380 44596 17382
rect 47582 21936 47638 21992
rect 51524 23418 51580 23420
rect 51604 23418 51660 23420
rect 51684 23418 51740 23420
rect 51764 23418 51820 23420
rect 51524 23366 51570 23418
rect 51570 23366 51580 23418
rect 51604 23366 51634 23418
rect 51634 23366 51646 23418
rect 51646 23366 51660 23418
rect 51684 23366 51698 23418
rect 51698 23366 51710 23418
rect 51710 23366 51740 23418
rect 51764 23366 51774 23418
rect 51774 23366 51820 23418
rect 51524 23364 51580 23366
rect 51604 23364 51660 23366
rect 51684 23364 51740 23366
rect 51764 23364 51820 23366
rect 44300 16346 44356 16348
rect 44380 16346 44436 16348
rect 44460 16346 44516 16348
rect 44540 16346 44596 16348
rect 44300 16294 44346 16346
rect 44346 16294 44356 16346
rect 44380 16294 44410 16346
rect 44410 16294 44422 16346
rect 44422 16294 44436 16346
rect 44460 16294 44474 16346
rect 44474 16294 44486 16346
rect 44486 16294 44516 16346
rect 44540 16294 44550 16346
rect 44550 16294 44596 16346
rect 44300 16292 44356 16294
rect 44380 16292 44436 16294
rect 44460 16292 44516 16294
rect 44540 16292 44596 16294
rect 44300 15258 44356 15260
rect 44380 15258 44436 15260
rect 44460 15258 44516 15260
rect 44540 15258 44596 15260
rect 44300 15206 44346 15258
rect 44346 15206 44356 15258
rect 44380 15206 44410 15258
rect 44410 15206 44422 15258
rect 44422 15206 44436 15258
rect 44460 15206 44474 15258
rect 44474 15206 44486 15258
rect 44486 15206 44516 15258
rect 44540 15206 44550 15258
rect 44550 15206 44596 15258
rect 44300 15204 44356 15206
rect 44380 15204 44436 15206
rect 44460 15204 44516 15206
rect 44540 15204 44596 15206
rect 45190 17176 45246 17232
rect 44300 14170 44356 14172
rect 44380 14170 44436 14172
rect 44460 14170 44516 14172
rect 44540 14170 44596 14172
rect 44300 14118 44346 14170
rect 44346 14118 44356 14170
rect 44380 14118 44410 14170
rect 44410 14118 44422 14170
rect 44422 14118 44436 14170
rect 44460 14118 44474 14170
rect 44474 14118 44486 14170
rect 44486 14118 44516 14170
rect 44540 14118 44550 14170
rect 44550 14118 44596 14170
rect 44300 14116 44356 14118
rect 44380 14116 44436 14118
rect 44460 14116 44516 14118
rect 44540 14116 44596 14118
rect 44300 13082 44356 13084
rect 44380 13082 44436 13084
rect 44460 13082 44516 13084
rect 44540 13082 44596 13084
rect 44300 13030 44346 13082
rect 44346 13030 44356 13082
rect 44380 13030 44410 13082
rect 44410 13030 44422 13082
rect 44422 13030 44436 13082
rect 44460 13030 44474 13082
rect 44474 13030 44486 13082
rect 44486 13030 44516 13082
rect 44540 13030 44550 13082
rect 44550 13030 44596 13082
rect 44300 13028 44356 13030
rect 44380 13028 44436 13030
rect 44460 13028 44516 13030
rect 44540 13028 44596 13030
rect 46846 18264 46902 18320
rect 44300 11994 44356 11996
rect 44380 11994 44436 11996
rect 44460 11994 44516 11996
rect 44540 11994 44596 11996
rect 44300 11942 44346 11994
rect 44346 11942 44356 11994
rect 44380 11942 44410 11994
rect 44410 11942 44422 11994
rect 44422 11942 44436 11994
rect 44460 11942 44474 11994
rect 44474 11942 44486 11994
rect 44486 11942 44516 11994
rect 44540 11942 44550 11994
rect 44550 11942 44596 11994
rect 44300 11940 44356 11942
rect 44380 11940 44436 11942
rect 44460 11940 44516 11942
rect 44540 11940 44596 11942
rect 44300 10906 44356 10908
rect 44380 10906 44436 10908
rect 44460 10906 44516 10908
rect 44540 10906 44596 10908
rect 44300 10854 44346 10906
rect 44346 10854 44356 10906
rect 44380 10854 44410 10906
rect 44410 10854 44422 10906
rect 44422 10854 44436 10906
rect 44460 10854 44474 10906
rect 44474 10854 44486 10906
rect 44486 10854 44516 10906
rect 44540 10854 44550 10906
rect 44550 10854 44596 10906
rect 44300 10852 44356 10854
rect 44380 10852 44436 10854
rect 44460 10852 44516 10854
rect 44540 10852 44596 10854
rect 44300 9818 44356 9820
rect 44380 9818 44436 9820
rect 44460 9818 44516 9820
rect 44540 9818 44596 9820
rect 44300 9766 44346 9818
rect 44346 9766 44356 9818
rect 44380 9766 44410 9818
rect 44410 9766 44422 9818
rect 44422 9766 44436 9818
rect 44460 9766 44474 9818
rect 44474 9766 44486 9818
rect 44486 9766 44516 9818
rect 44540 9766 44550 9818
rect 44550 9766 44596 9818
rect 44300 9764 44356 9766
rect 44380 9764 44436 9766
rect 44460 9764 44516 9766
rect 44540 9764 44596 9766
rect 44300 8730 44356 8732
rect 44380 8730 44436 8732
rect 44460 8730 44516 8732
rect 44540 8730 44596 8732
rect 44300 8678 44346 8730
rect 44346 8678 44356 8730
rect 44380 8678 44410 8730
rect 44410 8678 44422 8730
rect 44422 8678 44436 8730
rect 44460 8678 44474 8730
rect 44474 8678 44486 8730
rect 44486 8678 44516 8730
rect 44540 8678 44550 8730
rect 44550 8678 44596 8730
rect 44300 8676 44356 8678
rect 44380 8676 44436 8678
rect 44460 8676 44516 8678
rect 44540 8676 44596 8678
rect 43074 8236 43076 8256
rect 43076 8236 43128 8256
rect 43128 8236 43130 8256
rect 43074 8200 43130 8236
rect 42062 4528 42118 4584
rect 44300 7642 44356 7644
rect 44380 7642 44436 7644
rect 44460 7642 44516 7644
rect 44540 7642 44596 7644
rect 44300 7590 44346 7642
rect 44346 7590 44356 7642
rect 44380 7590 44410 7642
rect 44410 7590 44422 7642
rect 44422 7590 44436 7642
rect 44460 7590 44474 7642
rect 44474 7590 44486 7642
rect 44486 7590 44516 7642
rect 44540 7590 44550 7642
rect 44550 7590 44596 7642
rect 44300 7588 44356 7590
rect 44380 7588 44436 7590
rect 44460 7588 44516 7590
rect 44540 7588 44596 7590
rect 44822 8336 44878 8392
rect 51524 22330 51580 22332
rect 51604 22330 51660 22332
rect 51684 22330 51740 22332
rect 51764 22330 51820 22332
rect 51524 22278 51570 22330
rect 51570 22278 51580 22330
rect 51604 22278 51634 22330
rect 51634 22278 51646 22330
rect 51646 22278 51660 22330
rect 51684 22278 51698 22330
rect 51698 22278 51710 22330
rect 51710 22278 51740 22330
rect 51764 22278 51774 22330
rect 51774 22278 51820 22330
rect 51524 22276 51580 22278
rect 51604 22276 51660 22278
rect 51684 22276 51740 22278
rect 51764 22276 51820 22278
rect 48318 17720 48374 17776
rect 51524 21242 51580 21244
rect 51604 21242 51660 21244
rect 51684 21242 51740 21244
rect 51764 21242 51820 21244
rect 51524 21190 51570 21242
rect 51570 21190 51580 21242
rect 51604 21190 51634 21242
rect 51634 21190 51646 21242
rect 51646 21190 51660 21242
rect 51684 21190 51698 21242
rect 51698 21190 51710 21242
rect 51710 21190 51740 21242
rect 51764 21190 51774 21242
rect 51774 21190 51820 21242
rect 51524 21188 51580 21190
rect 51604 21188 51660 21190
rect 51684 21188 51740 21190
rect 51764 21188 51820 21190
rect 51524 20154 51580 20156
rect 51604 20154 51660 20156
rect 51684 20154 51740 20156
rect 51764 20154 51820 20156
rect 51524 20102 51570 20154
rect 51570 20102 51580 20154
rect 51604 20102 51634 20154
rect 51634 20102 51646 20154
rect 51646 20102 51660 20154
rect 51684 20102 51698 20154
rect 51698 20102 51710 20154
rect 51710 20102 51740 20154
rect 51764 20102 51774 20154
rect 51774 20102 51820 20154
rect 51524 20100 51580 20102
rect 51604 20100 51660 20102
rect 51684 20100 51740 20102
rect 51764 20100 51820 20102
rect 51524 19066 51580 19068
rect 51604 19066 51660 19068
rect 51684 19066 51740 19068
rect 51764 19066 51820 19068
rect 51524 19014 51570 19066
rect 51570 19014 51580 19066
rect 51604 19014 51634 19066
rect 51634 19014 51646 19066
rect 51646 19014 51660 19066
rect 51684 19014 51698 19066
rect 51698 19014 51710 19066
rect 51710 19014 51740 19066
rect 51764 19014 51774 19066
rect 51774 19014 51820 19066
rect 51524 19012 51580 19014
rect 51604 19012 51660 19014
rect 51684 19012 51740 19014
rect 51764 19012 51820 19014
rect 56598 21936 56654 21992
rect 46386 8200 46442 8256
rect 44300 6554 44356 6556
rect 44380 6554 44436 6556
rect 44460 6554 44516 6556
rect 44540 6554 44596 6556
rect 44300 6502 44346 6554
rect 44346 6502 44356 6554
rect 44380 6502 44410 6554
rect 44410 6502 44422 6554
rect 44422 6502 44436 6554
rect 44460 6502 44474 6554
rect 44474 6502 44486 6554
rect 44486 6502 44516 6554
rect 44540 6502 44550 6554
rect 44550 6502 44596 6554
rect 44300 6500 44356 6502
rect 44380 6500 44436 6502
rect 44460 6500 44516 6502
rect 44540 6500 44596 6502
rect 44300 5466 44356 5468
rect 44380 5466 44436 5468
rect 44460 5466 44516 5468
rect 44540 5466 44596 5468
rect 44300 5414 44346 5466
rect 44346 5414 44356 5466
rect 44380 5414 44410 5466
rect 44410 5414 44422 5466
rect 44422 5414 44436 5466
rect 44460 5414 44474 5466
rect 44474 5414 44486 5466
rect 44486 5414 44516 5466
rect 44540 5414 44550 5466
rect 44550 5414 44596 5466
rect 44300 5412 44356 5414
rect 44380 5412 44436 5414
rect 44460 5412 44516 5414
rect 44540 5412 44596 5414
rect 44300 4378 44356 4380
rect 44380 4378 44436 4380
rect 44460 4378 44516 4380
rect 44540 4378 44596 4380
rect 44300 4326 44346 4378
rect 44346 4326 44356 4378
rect 44380 4326 44410 4378
rect 44410 4326 44422 4378
rect 44422 4326 44436 4378
rect 44460 4326 44474 4378
rect 44474 4326 44486 4378
rect 44486 4326 44516 4378
rect 44540 4326 44550 4378
rect 44550 4326 44596 4378
rect 44300 4324 44356 4326
rect 44380 4324 44436 4326
rect 44460 4324 44516 4326
rect 44540 4324 44596 4326
rect 44300 3290 44356 3292
rect 44380 3290 44436 3292
rect 44460 3290 44516 3292
rect 44540 3290 44596 3292
rect 44300 3238 44346 3290
rect 44346 3238 44356 3290
rect 44380 3238 44410 3290
rect 44410 3238 44422 3290
rect 44422 3238 44436 3290
rect 44460 3238 44474 3290
rect 44474 3238 44486 3290
rect 44486 3238 44516 3290
rect 44540 3238 44550 3290
rect 44550 3238 44596 3290
rect 44300 3236 44356 3238
rect 44380 3236 44436 3238
rect 44460 3236 44516 3238
rect 44540 3236 44596 3238
rect 51524 17978 51580 17980
rect 51604 17978 51660 17980
rect 51684 17978 51740 17980
rect 51764 17978 51820 17980
rect 51524 17926 51570 17978
rect 51570 17926 51580 17978
rect 51604 17926 51634 17978
rect 51634 17926 51646 17978
rect 51646 17926 51660 17978
rect 51684 17926 51698 17978
rect 51698 17926 51710 17978
rect 51710 17926 51740 17978
rect 51764 17926 51774 17978
rect 51774 17926 51820 17978
rect 51524 17924 51580 17926
rect 51604 17924 51660 17926
rect 51684 17924 51740 17926
rect 51764 17924 51820 17926
rect 51906 17856 51962 17912
rect 51524 16890 51580 16892
rect 51604 16890 51660 16892
rect 51684 16890 51740 16892
rect 51764 16890 51820 16892
rect 51524 16838 51570 16890
rect 51570 16838 51580 16890
rect 51604 16838 51634 16890
rect 51634 16838 51646 16890
rect 51646 16838 51660 16890
rect 51684 16838 51698 16890
rect 51698 16838 51710 16890
rect 51710 16838 51740 16890
rect 51764 16838 51774 16890
rect 51774 16838 51820 16890
rect 51524 16836 51580 16838
rect 51604 16836 51660 16838
rect 51684 16836 51740 16838
rect 51764 16836 51820 16838
rect 51170 15952 51226 16008
rect 51524 15802 51580 15804
rect 51604 15802 51660 15804
rect 51684 15802 51740 15804
rect 51764 15802 51820 15804
rect 51524 15750 51570 15802
rect 51570 15750 51580 15802
rect 51604 15750 51634 15802
rect 51634 15750 51646 15802
rect 51646 15750 51660 15802
rect 51684 15750 51698 15802
rect 51698 15750 51710 15802
rect 51710 15750 51740 15802
rect 51764 15750 51774 15802
rect 51774 15750 51820 15802
rect 51524 15748 51580 15750
rect 51604 15748 51660 15750
rect 51684 15748 51740 15750
rect 51764 15748 51820 15750
rect 50618 15408 50674 15464
rect 50986 15408 51042 15464
rect 51524 14714 51580 14716
rect 51604 14714 51660 14716
rect 51684 14714 51740 14716
rect 51764 14714 51820 14716
rect 51524 14662 51570 14714
rect 51570 14662 51580 14714
rect 51604 14662 51634 14714
rect 51634 14662 51646 14714
rect 51646 14662 51660 14714
rect 51684 14662 51698 14714
rect 51698 14662 51710 14714
rect 51710 14662 51740 14714
rect 51764 14662 51774 14714
rect 51774 14662 51820 14714
rect 51524 14660 51580 14662
rect 51604 14660 51660 14662
rect 51684 14660 51740 14662
rect 51764 14660 51820 14662
rect 51524 13626 51580 13628
rect 51604 13626 51660 13628
rect 51684 13626 51740 13628
rect 51764 13626 51820 13628
rect 51524 13574 51570 13626
rect 51570 13574 51580 13626
rect 51604 13574 51634 13626
rect 51634 13574 51646 13626
rect 51646 13574 51660 13626
rect 51684 13574 51698 13626
rect 51698 13574 51710 13626
rect 51710 13574 51740 13626
rect 51764 13574 51774 13626
rect 51774 13574 51820 13626
rect 51524 13572 51580 13574
rect 51604 13572 51660 13574
rect 51684 13572 51740 13574
rect 51764 13572 51820 13574
rect 51524 12538 51580 12540
rect 51604 12538 51660 12540
rect 51684 12538 51740 12540
rect 51764 12538 51820 12540
rect 51524 12486 51570 12538
rect 51570 12486 51580 12538
rect 51604 12486 51634 12538
rect 51634 12486 51646 12538
rect 51646 12486 51660 12538
rect 51684 12486 51698 12538
rect 51698 12486 51710 12538
rect 51710 12486 51740 12538
rect 51764 12486 51774 12538
rect 51774 12486 51820 12538
rect 51524 12484 51580 12486
rect 51604 12484 51660 12486
rect 51684 12484 51740 12486
rect 51764 12484 51820 12486
rect 52826 15408 52882 15464
rect 53838 17856 53894 17912
rect 57242 17060 57298 17096
rect 57242 17040 57244 17060
rect 57244 17040 57296 17060
rect 57296 17040 57298 17060
rect 57058 15988 57060 16008
rect 57060 15988 57112 16008
rect 57112 15988 57114 16008
rect 57058 15952 57114 15988
rect 51524 11450 51580 11452
rect 51604 11450 51660 11452
rect 51684 11450 51740 11452
rect 51764 11450 51820 11452
rect 51524 11398 51570 11450
rect 51570 11398 51580 11450
rect 51604 11398 51634 11450
rect 51634 11398 51646 11450
rect 51646 11398 51660 11450
rect 51684 11398 51698 11450
rect 51698 11398 51710 11450
rect 51710 11398 51740 11450
rect 51764 11398 51774 11450
rect 51774 11398 51820 11450
rect 51524 11396 51580 11398
rect 51604 11396 51660 11398
rect 51684 11396 51740 11398
rect 51764 11396 51820 11398
rect 51524 10362 51580 10364
rect 51604 10362 51660 10364
rect 51684 10362 51740 10364
rect 51764 10362 51820 10364
rect 51524 10310 51570 10362
rect 51570 10310 51580 10362
rect 51604 10310 51634 10362
rect 51634 10310 51646 10362
rect 51646 10310 51660 10362
rect 51684 10310 51698 10362
rect 51698 10310 51710 10362
rect 51710 10310 51740 10362
rect 51764 10310 51774 10362
rect 51774 10310 51820 10362
rect 51524 10308 51580 10310
rect 51604 10308 51660 10310
rect 51684 10308 51740 10310
rect 51764 10308 51820 10310
rect 51524 9274 51580 9276
rect 51604 9274 51660 9276
rect 51684 9274 51740 9276
rect 51764 9274 51820 9276
rect 51524 9222 51570 9274
rect 51570 9222 51580 9274
rect 51604 9222 51634 9274
rect 51634 9222 51646 9274
rect 51646 9222 51660 9274
rect 51684 9222 51698 9274
rect 51698 9222 51710 9274
rect 51710 9222 51740 9274
rect 51764 9222 51774 9274
rect 51774 9222 51820 9274
rect 51524 9220 51580 9222
rect 51604 9220 51660 9222
rect 51684 9220 51740 9222
rect 51764 9220 51820 9222
rect 55402 9560 55458 9616
rect 55586 8880 55642 8936
rect 58070 33380 58126 33416
rect 58070 33360 58072 33380
rect 58072 33360 58124 33380
rect 58124 33360 58126 33380
rect 58070 27920 58126 27976
rect 57886 23160 57942 23216
rect 57794 17720 57850 17776
rect 57610 11056 57666 11112
rect 51524 8186 51580 8188
rect 51604 8186 51660 8188
rect 51684 8186 51740 8188
rect 51764 8186 51820 8188
rect 51524 8134 51570 8186
rect 51570 8134 51580 8186
rect 51604 8134 51634 8186
rect 51634 8134 51646 8186
rect 51646 8134 51660 8186
rect 51684 8134 51698 8186
rect 51698 8134 51710 8186
rect 51710 8134 51740 8186
rect 51764 8134 51774 8186
rect 51774 8134 51820 8186
rect 51524 8132 51580 8134
rect 51604 8132 51660 8134
rect 51684 8132 51740 8134
rect 51764 8132 51820 8134
rect 51524 7098 51580 7100
rect 51604 7098 51660 7100
rect 51684 7098 51740 7100
rect 51764 7098 51820 7100
rect 51524 7046 51570 7098
rect 51570 7046 51580 7098
rect 51604 7046 51634 7098
rect 51634 7046 51646 7098
rect 51646 7046 51660 7098
rect 51684 7046 51698 7098
rect 51698 7046 51710 7098
rect 51710 7046 51740 7098
rect 51764 7046 51774 7098
rect 51774 7046 51820 7098
rect 51524 7044 51580 7046
rect 51604 7044 51660 7046
rect 51684 7044 51740 7046
rect 51764 7044 51820 7046
rect 51524 6010 51580 6012
rect 51604 6010 51660 6012
rect 51684 6010 51740 6012
rect 51764 6010 51820 6012
rect 51524 5958 51570 6010
rect 51570 5958 51580 6010
rect 51604 5958 51634 6010
rect 51634 5958 51646 6010
rect 51646 5958 51660 6010
rect 51684 5958 51698 6010
rect 51698 5958 51710 6010
rect 51710 5958 51740 6010
rect 51764 5958 51774 6010
rect 51774 5958 51820 6010
rect 51524 5956 51580 5958
rect 51604 5956 51660 5958
rect 51684 5956 51740 5958
rect 51764 5956 51820 5958
rect 51524 4922 51580 4924
rect 51604 4922 51660 4924
rect 51684 4922 51740 4924
rect 51764 4922 51820 4924
rect 51524 4870 51570 4922
rect 51570 4870 51580 4922
rect 51604 4870 51634 4922
rect 51634 4870 51646 4922
rect 51646 4870 51660 4922
rect 51684 4870 51698 4922
rect 51698 4870 51710 4922
rect 51710 4870 51740 4922
rect 51764 4870 51774 4922
rect 51774 4870 51820 4922
rect 51524 4868 51580 4870
rect 51604 4868 51660 4870
rect 51684 4868 51740 4870
rect 51764 4868 51820 4870
rect 51524 3834 51580 3836
rect 51604 3834 51660 3836
rect 51684 3834 51740 3836
rect 51764 3834 51820 3836
rect 51524 3782 51570 3834
rect 51570 3782 51580 3834
rect 51604 3782 51634 3834
rect 51634 3782 51646 3834
rect 51646 3782 51660 3834
rect 51684 3782 51698 3834
rect 51698 3782 51710 3834
rect 51710 3782 51740 3834
rect 51764 3782 51774 3834
rect 51774 3782 51820 3834
rect 51524 3780 51580 3782
rect 51604 3780 51660 3782
rect 51684 3780 51740 3782
rect 51764 3780 51820 3782
rect 51524 2746 51580 2748
rect 51604 2746 51660 2748
rect 51684 2746 51740 2748
rect 51764 2746 51820 2748
rect 51524 2694 51570 2746
rect 51570 2694 51580 2746
rect 51604 2694 51634 2746
rect 51634 2694 51646 2746
rect 51646 2694 51660 2746
rect 51684 2694 51698 2746
rect 51698 2694 51710 2746
rect 51710 2694 51740 2746
rect 51764 2694 51774 2746
rect 51774 2694 51820 2746
rect 51524 2692 51580 2694
rect 51604 2692 51660 2694
rect 51684 2692 51740 2694
rect 51764 2692 51820 2694
rect 15404 2202 15460 2204
rect 15484 2202 15540 2204
rect 15564 2202 15620 2204
rect 15644 2202 15700 2204
rect 15404 2150 15450 2202
rect 15450 2150 15460 2202
rect 15484 2150 15514 2202
rect 15514 2150 15526 2202
rect 15526 2150 15540 2202
rect 15564 2150 15578 2202
rect 15578 2150 15590 2202
rect 15590 2150 15620 2202
rect 15644 2150 15654 2202
rect 15654 2150 15700 2202
rect 15404 2148 15460 2150
rect 15484 2148 15540 2150
rect 15564 2148 15620 2150
rect 15644 2148 15700 2150
rect 29852 2202 29908 2204
rect 29932 2202 29988 2204
rect 30012 2202 30068 2204
rect 30092 2202 30148 2204
rect 29852 2150 29898 2202
rect 29898 2150 29908 2202
rect 29932 2150 29962 2202
rect 29962 2150 29974 2202
rect 29974 2150 29988 2202
rect 30012 2150 30026 2202
rect 30026 2150 30038 2202
rect 30038 2150 30068 2202
rect 30092 2150 30102 2202
rect 30102 2150 30148 2202
rect 29852 2148 29908 2150
rect 29932 2148 29988 2150
rect 30012 2148 30068 2150
rect 30092 2148 30148 2150
rect 58070 12980 58126 13016
rect 58070 12960 58072 12980
rect 58072 12960 58124 12980
rect 58124 12960 58126 12980
rect 58070 7520 58126 7576
rect 58070 2796 58072 2816
rect 58072 2796 58124 2816
rect 58124 2796 58126 2816
rect 58070 2760 58126 2796
rect 44300 2202 44356 2204
rect 44380 2202 44436 2204
rect 44460 2202 44516 2204
rect 44540 2202 44596 2204
rect 44300 2150 44346 2202
rect 44346 2150 44356 2202
rect 44380 2150 44410 2202
rect 44410 2150 44422 2202
rect 44422 2150 44436 2202
rect 44460 2150 44474 2202
rect 44474 2150 44486 2202
rect 44486 2150 44516 2202
rect 44540 2150 44550 2202
rect 44550 2150 44596 2202
rect 44300 2148 44356 2150
rect 44380 2148 44436 2150
rect 44460 2148 44516 2150
rect 44540 2148 44596 2150
<< metal3 >>
rect 0 35458 800 35488
rect 1485 35458 1551 35461
rect 0 35456 1551 35458
rect 0 35400 1490 35456
rect 1546 35400 1551 35456
rect 0 35398 1551 35400
rect 0 35368 800 35398
rect 1485 35395 1551 35398
rect 15394 33760 15710 33761
rect 15394 33696 15400 33760
rect 15464 33696 15480 33760
rect 15544 33696 15560 33760
rect 15624 33696 15640 33760
rect 15704 33696 15710 33760
rect 15394 33695 15710 33696
rect 29842 33760 30158 33761
rect 29842 33696 29848 33760
rect 29912 33696 29928 33760
rect 29992 33696 30008 33760
rect 30072 33696 30088 33760
rect 30152 33696 30158 33760
rect 29842 33695 30158 33696
rect 44290 33760 44606 33761
rect 44290 33696 44296 33760
rect 44360 33696 44376 33760
rect 44440 33696 44456 33760
rect 44520 33696 44536 33760
rect 44600 33696 44606 33760
rect 44290 33695 44606 33696
rect 58065 33418 58131 33421
rect 59200 33418 60000 33448
rect 58065 33416 60000 33418
rect 58065 33360 58070 33416
rect 58126 33360 60000 33416
rect 58065 33358 60000 33360
rect 58065 33355 58131 33358
rect 59200 33328 60000 33358
rect 8170 33216 8486 33217
rect 8170 33152 8176 33216
rect 8240 33152 8256 33216
rect 8320 33152 8336 33216
rect 8400 33152 8416 33216
rect 8480 33152 8486 33216
rect 8170 33151 8486 33152
rect 22618 33216 22934 33217
rect 22618 33152 22624 33216
rect 22688 33152 22704 33216
rect 22768 33152 22784 33216
rect 22848 33152 22864 33216
rect 22928 33152 22934 33216
rect 22618 33151 22934 33152
rect 37066 33216 37382 33217
rect 37066 33152 37072 33216
rect 37136 33152 37152 33216
rect 37216 33152 37232 33216
rect 37296 33152 37312 33216
rect 37376 33152 37382 33216
rect 37066 33151 37382 33152
rect 51514 33216 51830 33217
rect 51514 33152 51520 33216
rect 51584 33152 51600 33216
rect 51664 33152 51680 33216
rect 51744 33152 51760 33216
rect 51824 33152 51830 33216
rect 51514 33151 51830 33152
rect 15394 32672 15710 32673
rect 15394 32608 15400 32672
rect 15464 32608 15480 32672
rect 15544 32608 15560 32672
rect 15624 32608 15640 32672
rect 15704 32608 15710 32672
rect 15394 32607 15710 32608
rect 29842 32672 30158 32673
rect 29842 32608 29848 32672
rect 29912 32608 29928 32672
rect 29992 32608 30008 32672
rect 30072 32608 30088 32672
rect 30152 32608 30158 32672
rect 29842 32607 30158 32608
rect 44290 32672 44606 32673
rect 44290 32608 44296 32672
rect 44360 32608 44376 32672
rect 44440 32608 44456 32672
rect 44520 32608 44536 32672
rect 44600 32608 44606 32672
rect 44290 32607 44606 32608
rect 8170 32128 8486 32129
rect 8170 32064 8176 32128
rect 8240 32064 8256 32128
rect 8320 32064 8336 32128
rect 8400 32064 8416 32128
rect 8480 32064 8486 32128
rect 8170 32063 8486 32064
rect 22618 32128 22934 32129
rect 22618 32064 22624 32128
rect 22688 32064 22704 32128
rect 22768 32064 22784 32128
rect 22848 32064 22864 32128
rect 22928 32064 22934 32128
rect 22618 32063 22934 32064
rect 37066 32128 37382 32129
rect 37066 32064 37072 32128
rect 37136 32064 37152 32128
rect 37216 32064 37232 32128
rect 37296 32064 37312 32128
rect 37376 32064 37382 32128
rect 37066 32063 37382 32064
rect 51514 32128 51830 32129
rect 51514 32064 51520 32128
rect 51584 32064 51600 32128
rect 51664 32064 51680 32128
rect 51744 32064 51760 32128
rect 51824 32064 51830 32128
rect 51514 32063 51830 32064
rect 15394 31584 15710 31585
rect 15394 31520 15400 31584
rect 15464 31520 15480 31584
rect 15544 31520 15560 31584
rect 15624 31520 15640 31584
rect 15704 31520 15710 31584
rect 15394 31519 15710 31520
rect 29842 31584 30158 31585
rect 29842 31520 29848 31584
rect 29912 31520 29928 31584
rect 29992 31520 30008 31584
rect 30072 31520 30088 31584
rect 30152 31520 30158 31584
rect 29842 31519 30158 31520
rect 44290 31584 44606 31585
rect 44290 31520 44296 31584
rect 44360 31520 44376 31584
rect 44440 31520 44456 31584
rect 44520 31520 44536 31584
rect 44600 31520 44606 31584
rect 44290 31519 44606 31520
rect 8170 31040 8486 31041
rect 8170 30976 8176 31040
rect 8240 30976 8256 31040
rect 8320 30976 8336 31040
rect 8400 30976 8416 31040
rect 8480 30976 8486 31040
rect 8170 30975 8486 30976
rect 22618 31040 22934 31041
rect 22618 30976 22624 31040
rect 22688 30976 22704 31040
rect 22768 30976 22784 31040
rect 22848 30976 22864 31040
rect 22928 30976 22934 31040
rect 22618 30975 22934 30976
rect 37066 31040 37382 31041
rect 37066 30976 37072 31040
rect 37136 30976 37152 31040
rect 37216 30976 37232 31040
rect 37296 30976 37312 31040
rect 37376 30976 37382 31040
rect 37066 30975 37382 30976
rect 51514 31040 51830 31041
rect 51514 30976 51520 31040
rect 51584 30976 51600 31040
rect 51664 30976 51680 31040
rect 51744 30976 51760 31040
rect 51824 30976 51830 31040
rect 51514 30975 51830 30976
rect 0 30698 800 30728
rect 1485 30698 1551 30701
rect 0 30696 1551 30698
rect 0 30640 1490 30696
rect 1546 30640 1551 30696
rect 0 30638 1551 30640
rect 0 30608 800 30638
rect 1485 30635 1551 30638
rect 15394 30496 15710 30497
rect 15394 30432 15400 30496
rect 15464 30432 15480 30496
rect 15544 30432 15560 30496
rect 15624 30432 15640 30496
rect 15704 30432 15710 30496
rect 15394 30431 15710 30432
rect 29842 30496 30158 30497
rect 29842 30432 29848 30496
rect 29912 30432 29928 30496
rect 29992 30432 30008 30496
rect 30072 30432 30088 30496
rect 30152 30432 30158 30496
rect 29842 30431 30158 30432
rect 44290 30496 44606 30497
rect 44290 30432 44296 30496
rect 44360 30432 44376 30496
rect 44440 30432 44456 30496
rect 44520 30432 44536 30496
rect 44600 30432 44606 30496
rect 44290 30431 44606 30432
rect 8170 29952 8486 29953
rect 8170 29888 8176 29952
rect 8240 29888 8256 29952
rect 8320 29888 8336 29952
rect 8400 29888 8416 29952
rect 8480 29888 8486 29952
rect 8170 29887 8486 29888
rect 22618 29952 22934 29953
rect 22618 29888 22624 29952
rect 22688 29888 22704 29952
rect 22768 29888 22784 29952
rect 22848 29888 22864 29952
rect 22928 29888 22934 29952
rect 22618 29887 22934 29888
rect 37066 29952 37382 29953
rect 37066 29888 37072 29952
rect 37136 29888 37152 29952
rect 37216 29888 37232 29952
rect 37296 29888 37312 29952
rect 37376 29888 37382 29952
rect 37066 29887 37382 29888
rect 51514 29952 51830 29953
rect 51514 29888 51520 29952
rect 51584 29888 51600 29952
rect 51664 29888 51680 29952
rect 51744 29888 51760 29952
rect 51824 29888 51830 29952
rect 51514 29887 51830 29888
rect 15394 29408 15710 29409
rect 15394 29344 15400 29408
rect 15464 29344 15480 29408
rect 15544 29344 15560 29408
rect 15624 29344 15640 29408
rect 15704 29344 15710 29408
rect 15394 29343 15710 29344
rect 29842 29408 30158 29409
rect 29842 29344 29848 29408
rect 29912 29344 29928 29408
rect 29992 29344 30008 29408
rect 30072 29344 30088 29408
rect 30152 29344 30158 29408
rect 29842 29343 30158 29344
rect 44290 29408 44606 29409
rect 44290 29344 44296 29408
rect 44360 29344 44376 29408
rect 44440 29344 44456 29408
rect 44520 29344 44536 29408
rect 44600 29344 44606 29408
rect 44290 29343 44606 29344
rect 8170 28864 8486 28865
rect 8170 28800 8176 28864
rect 8240 28800 8256 28864
rect 8320 28800 8336 28864
rect 8400 28800 8416 28864
rect 8480 28800 8486 28864
rect 8170 28799 8486 28800
rect 22618 28864 22934 28865
rect 22618 28800 22624 28864
rect 22688 28800 22704 28864
rect 22768 28800 22784 28864
rect 22848 28800 22864 28864
rect 22928 28800 22934 28864
rect 22618 28799 22934 28800
rect 37066 28864 37382 28865
rect 37066 28800 37072 28864
rect 37136 28800 37152 28864
rect 37216 28800 37232 28864
rect 37296 28800 37312 28864
rect 37376 28800 37382 28864
rect 37066 28799 37382 28800
rect 51514 28864 51830 28865
rect 51514 28800 51520 28864
rect 51584 28800 51600 28864
rect 51664 28800 51680 28864
rect 51744 28800 51760 28864
rect 51824 28800 51830 28864
rect 51514 28799 51830 28800
rect 15394 28320 15710 28321
rect 15394 28256 15400 28320
rect 15464 28256 15480 28320
rect 15544 28256 15560 28320
rect 15624 28256 15640 28320
rect 15704 28256 15710 28320
rect 15394 28255 15710 28256
rect 29842 28320 30158 28321
rect 29842 28256 29848 28320
rect 29912 28256 29928 28320
rect 29992 28256 30008 28320
rect 30072 28256 30088 28320
rect 30152 28256 30158 28320
rect 29842 28255 30158 28256
rect 44290 28320 44606 28321
rect 44290 28256 44296 28320
rect 44360 28256 44376 28320
rect 44440 28256 44456 28320
rect 44520 28256 44536 28320
rect 44600 28256 44606 28320
rect 44290 28255 44606 28256
rect 4245 27978 4311 27981
rect 9029 27978 9095 27981
rect 4245 27976 9095 27978
rect 4245 27920 4250 27976
rect 4306 27920 9034 27976
rect 9090 27920 9095 27976
rect 4245 27918 9095 27920
rect 4245 27915 4311 27918
rect 9029 27915 9095 27918
rect 58065 27978 58131 27981
rect 59200 27978 60000 28008
rect 58065 27976 60000 27978
rect 58065 27920 58070 27976
rect 58126 27920 60000 27976
rect 58065 27918 60000 27920
rect 58065 27915 58131 27918
rect 59200 27888 60000 27918
rect 8170 27776 8486 27777
rect 8170 27712 8176 27776
rect 8240 27712 8256 27776
rect 8320 27712 8336 27776
rect 8400 27712 8416 27776
rect 8480 27712 8486 27776
rect 8170 27711 8486 27712
rect 22618 27776 22934 27777
rect 22618 27712 22624 27776
rect 22688 27712 22704 27776
rect 22768 27712 22784 27776
rect 22848 27712 22864 27776
rect 22928 27712 22934 27776
rect 22618 27711 22934 27712
rect 37066 27776 37382 27777
rect 37066 27712 37072 27776
rect 37136 27712 37152 27776
rect 37216 27712 37232 27776
rect 37296 27712 37312 27776
rect 37376 27712 37382 27776
rect 37066 27711 37382 27712
rect 51514 27776 51830 27777
rect 51514 27712 51520 27776
rect 51584 27712 51600 27776
rect 51664 27712 51680 27776
rect 51744 27712 51760 27776
rect 51824 27712 51830 27776
rect 51514 27711 51830 27712
rect 15394 27232 15710 27233
rect 15394 27168 15400 27232
rect 15464 27168 15480 27232
rect 15544 27168 15560 27232
rect 15624 27168 15640 27232
rect 15704 27168 15710 27232
rect 15394 27167 15710 27168
rect 29842 27232 30158 27233
rect 29842 27168 29848 27232
rect 29912 27168 29928 27232
rect 29992 27168 30008 27232
rect 30072 27168 30088 27232
rect 30152 27168 30158 27232
rect 29842 27167 30158 27168
rect 44290 27232 44606 27233
rect 44290 27168 44296 27232
rect 44360 27168 44376 27232
rect 44440 27168 44456 27232
rect 44520 27168 44536 27232
rect 44600 27168 44606 27232
rect 44290 27167 44606 27168
rect 8170 26688 8486 26689
rect 8170 26624 8176 26688
rect 8240 26624 8256 26688
rect 8320 26624 8336 26688
rect 8400 26624 8416 26688
rect 8480 26624 8486 26688
rect 8170 26623 8486 26624
rect 22618 26688 22934 26689
rect 22618 26624 22624 26688
rect 22688 26624 22704 26688
rect 22768 26624 22784 26688
rect 22848 26624 22864 26688
rect 22928 26624 22934 26688
rect 22618 26623 22934 26624
rect 37066 26688 37382 26689
rect 37066 26624 37072 26688
rect 37136 26624 37152 26688
rect 37216 26624 37232 26688
rect 37296 26624 37312 26688
rect 37376 26624 37382 26688
rect 37066 26623 37382 26624
rect 51514 26688 51830 26689
rect 51514 26624 51520 26688
rect 51584 26624 51600 26688
rect 51664 26624 51680 26688
rect 51744 26624 51760 26688
rect 51824 26624 51830 26688
rect 51514 26623 51830 26624
rect 15394 26144 15710 26145
rect 15394 26080 15400 26144
rect 15464 26080 15480 26144
rect 15544 26080 15560 26144
rect 15624 26080 15640 26144
rect 15704 26080 15710 26144
rect 15394 26079 15710 26080
rect 29842 26144 30158 26145
rect 29842 26080 29848 26144
rect 29912 26080 29928 26144
rect 29992 26080 30008 26144
rect 30072 26080 30088 26144
rect 30152 26080 30158 26144
rect 29842 26079 30158 26080
rect 44290 26144 44606 26145
rect 44290 26080 44296 26144
rect 44360 26080 44376 26144
rect 44440 26080 44456 26144
rect 44520 26080 44536 26144
rect 44600 26080 44606 26144
rect 44290 26079 44606 26080
rect 8170 25600 8486 25601
rect 8170 25536 8176 25600
rect 8240 25536 8256 25600
rect 8320 25536 8336 25600
rect 8400 25536 8416 25600
rect 8480 25536 8486 25600
rect 8170 25535 8486 25536
rect 22618 25600 22934 25601
rect 22618 25536 22624 25600
rect 22688 25536 22704 25600
rect 22768 25536 22784 25600
rect 22848 25536 22864 25600
rect 22928 25536 22934 25600
rect 22618 25535 22934 25536
rect 37066 25600 37382 25601
rect 37066 25536 37072 25600
rect 37136 25536 37152 25600
rect 37216 25536 37232 25600
rect 37296 25536 37312 25600
rect 37376 25536 37382 25600
rect 37066 25535 37382 25536
rect 51514 25600 51830 25601
rect 51514 25536 51520 25600
rect 51584 25536 51600 25600
rect 51664 25536 51680 25600
rect 51744 25536 51760 25600
rect 51824 25536 51830 25600
rect 51514 25535 51830 25536
rect 12617 25394 12683 25397
rect 26325 25394 26391 25397
rect 12617 25392 26391 25394
rect 12617 25336 12622 25392
rect 12678 25336 26330 25392
rect 26386 25336 26391 25392
rect 12617 25334 26391 25336
rect 12617 25331 12683 25334
rect 26325 25331 26391 25334
rect 0 25258 800 25288
rect 1485 25258 1551 25261
rect 0 25256 1551 25258
rect 0 25200 1490 25256
rect 1546 25200 1551 25256
rect 0 25198 1551 25200
rect 0 25168 800 25198
rect 1485 25195 1551 25198
rect 17401 25258 17467 25261
rect 18321 25258 18387 25261
rect 17401 25256 18387 25258
rect 17401 25200 17406 25256
rect 17462 25200 18326 25256
rect 18382 25200 18387 25256
rect 17401 25198 18387 25200
rect 17401 25195 17467 25198
rect 18321 25195 18387 25198
rect 15394 25056 15710 25057
rect 15394 24992 15400 25056
rect 15464 24992 15480 25056
rect 15544 24992 15560 25056
rect 15624 24992 15640 25056
rect 15704 24992 15710 25056
rect 15394 24991 15710 24992
rect 29842 25056 30158 25057
rect 29842 24992 29848 25056
rect 29912 24992 29928 25056
rect 29992 24992 30008 25056
rect 30072 24992 30088 25056
rect 30152 24992 30158 25056
rect 29842 24991 30158 24992
rect 44290 25056 44606 25057
rect 44290 24992 44296 25056
rect 44360 24992 44376 25056
rect 44440 24992 44456 25056
rect 44520 24992 44536 25056
rect 44600 24992 44606 25056
rect 44290 24991 44606 24992
rect 2405 24850 2471 24853
rect 24485 24850 24551 24853
rect 2405 24848 24551 24850
rect 2405 24792 2410 24848
rect 2466 24792 24490 24848
rect 24546 24792 24551 24848
rect 2405 24790 24551 24792
rect 2405 24787 2471 24790
rect 24485 24787 24551 24790
rect 20805 24714 20871 24717
rect 37365 24714 37431 24717
rect 20805 24712 37431 24714
rect 20805 24656 20810 24712
rect 20866 24656 37370 24712
rect 37426 24656 37431 24712
rect 20805 24654 37431 24656
rect 20805 24651 20871 24654
rect 37365 24651 37431 24654
rect 8170 24512 8486 24513
rect 8170 24448 8176 24512
rect 8240 24448 8256 24512
rect 8320 24448 8336 24512
rect 8400 24448 8416 24512
rect 8480 24448 8486 24512
rect 8170 24447 8486 24448
rect 22618 24512 22934 24513
rect 22618 24448 22624 24512
rect 22688 24448 22704 24512
rect 22768 24448 22784 24512
rect 22848 24448 22864 24512
rect 22928 24448 22934 24512
rect 22618 24447 22934 24448
rect 37066 24512 37382 24513
rect 37066 24448 37072 24512
rect 37136 24448 37152 24512
rect 37216 24448 37232 24512
rect 37296 24448 37312 24512
rect 37376 24448 37382 24512
rect 37066 24447 37382 24448
rect 51514 24512 51830 24513
rect 51514 24448 51520 24512
rect 51584 24448 51600 24512
rect 51664 24448 51680 24512
rect 51744 24448 51760 24512
rect 51824 24448 51830 24512
rect 51514 24447 51830 24448
rect 8109 24306 8175 24309
rect 20529 24306 20595 24309
rect 8109 24304 20595 24306
rect 8109 24248 8114 24304
rect 8170 24248 20534 24304
rect 20590 24248 20595 24304
rect 8109 24246 20595 24248
rect 8109 24243 8175 24246
rect 20529 24243 20595 24246
rect 13629 24170 13695 24173
rect 21357 24170 21423 24173
rect 27429 24170 27495 24173
rect 13629 24168 27495 24170
rect 13629 24112 13634 24168
rect 13690 24112 21362 24168
rect 21418 24112 27434 24168
rect 27490 24112 27495 24168
rect 13629 24110 27495 24112
rect 13629 24107 13695 24110
rect 21357 24107 21423 24110
rect 27429 24107 27495 24110
rect 15394 23968 15710 23969
rect 15394 23904 15400 23968
rect 15464 23904 15480 23968
rect 15544 23904 15560 23968
rect 15624 23904 15640 23968
rect 15704 23904 15710 23968
rect 15394 23903 15710 23904
rect 29842 23968 30158 23969
rect 29842 23904 29848 23968
rect 29912 23904 29928 23968
rect 29992 23904 30008 23968
rect 30072 23904 30088 23968
rect 30152 23904 30158 23968
rect 29842 23903 30158 23904
rect 44290 23968 44606 23969
rect 44290 23904 44296 23968
rect 44360 23904 44376 23968
rect 44440 23904 44456 23968
rect 44520 23904 44536 23968
rect 44600 23904 44606 23968
rect 44290 23903 44606 23904
rect 19885 23762 19951 23765
rect 33593 23762 33659 23765
rect 19885 23760 33659 23762
rect 19885 23704 19890 23760
rect 19946 23704 33598 23760
rect 33654 23704 33659 23760
rect 19885 23702 33659 23704
rect 19885 23699 19951 23702
rect 33593 23699 33659 23702
rect 5809 23626 5875 23629
rect 21081 23626 21147 23629
rect 5809 23624 21147 23626
rect 5809 23568 5814 23624
rect 5870 23568 21086 23624
rect 21142 23568 21147 23624
rect 5809 23566 21147 23568
rect 5809 23563 5875 23566
rect 21081 23563 21147 23566
rect 8170 23424 8486 23425
rect 8170 23360 8176 23424
rect 8240 23360 8256 23424
rect 8320 23360 8336 23424
rect 8400 23360 8416 23424
rect 8480 23360 8486 23424
rect 8170 23359 8486 23360
rect 22618 23424 22934 23425
rect 22618 23360 22624 23424
rect 22688 23360 22704 23424
rect 22768 23360 22784 23424
rect 22848 23360 22864 23424
rect 22928 23360 22934 23424
rect 22618 23359 22934 23360
rect 37066 23424 37382 23425
rect 37066 23360 37072 23424
rect 37136 23360 37152 23424
rect 37216 23360 37232 23424
rect 37296 23360 37312 23424
rect 37376 23360 37382 23424
rect 37066 23359 37382 23360
rect 51514 23424 51830 23425
rect 51514 23360 51520 23424
rect 51584 23360 51600 23424
rect 51664 23360 51680 23424
rect 51744 23360 51760 23424
rect 51824 23360 51830 23424
rect 51514 23359 51830 23360
rect 2037 23218 2103 23221
rect 18413 23218 18479 23221
rect 2037 23216 18479 23218
rect 2037 23160 2042 23216
rect 2098 23160 18418 23216
rect 18474 23160 18479 23216
rect 2037 23158 18479 23160
rect 2037 23155 2103 23158
rect 18413 23155 18479 23158
rect 20713 23218 20779 23221
rect 25497 23218 25563 23221
rect 20713 23216 25563 23218
rect 20713 23160 20718 23216
rect 20774 23160 25502 23216
rect 25558 23160 25563 23216
rect 20713 23158 25563 23160
rect 20713 23155 20779 23158
rect 25497 23155 25563 23158
rect 57881 23218 57947 23221
rect 59200 23218 60000 23248
rect 57881 23216 60000 23218
rect 57881 23160 57886 23216
rect 57942 23160 60000 23216
rect 57881 23158 60000 23160
rect 57881 23155 57947 23158
rect 59200 23128 60000 23158
rect 4889 23082 4955 23085
rect 18045 23082 18111 23085
rect 4889 23080 18111 23082
rect 4889 23024 4894 23080
rect 4950 23024 18050 23080
rect 18106 23024 18111 23080
rect 4889 23022 18111 23024
rect 4889 23019 4955 23022
rect 18045 23019 18111 23022
rect 24485 23082 24551 23085
rect 25221 23082 25287 23085
rect 26877 23082 26943 23085
rect 24485 23080 26943 23082
rect 24485 23024 24490 23080
rect 24546 23024 25226 23080
rect 25282 23024 26882 23080
rect 26938 23024 26943 23080
rect 24485 23022 26943 23024
rect 24485 23019 24551 23022
rect 25221 23019 25287 23022
rect 26877 23019 26943 23022
rect 15394 22880 15710 22881
rect 15394 22816 15400 22880
rect 15464 22816 15480 22880
rect 15544 22816 15560 22880
rect 15624 22816 15640 22880
rect 15704 22816 15710 22880
rect 15394 22815 15710 22816
rect 29842 22880 30158 22881
rect 29842 22816 29848 22880
rect 29912 22816 29928 22880
rect 29992 22816 30008 22880
rect 30072 22816 30088 22880
rect 30152 22816 30158 22880
rect 29842 22815 30158 22816
rect 44290 22880 44606 22881
rect 44290 22816 44296 22880
rect 44360 22816 44376 22880
rect 44440 22816 44456 22880
rect 44520 22816 44536 22880
rect 44600 22816 44606 22880
rect 44290 22815 44606 22816
rect 7373 22674 7439 22677
rect 17217 22674 17283 22677
rect 7373 22672 17283 22674
rect 7373 22616 7378 22672
rect 7434 22616 17222 22672
rect 17278 22616 17283 22672
rect 7373 22614 17283 22616
rect 7373 22611 7439 22614
rect 17217 22611 17283 22614
rect 18413 22538 18479 22541
rect 32949 22538 33015 22541
rect 18413 22536 33015 22538
rect 18413 22480 18418 22536
rect 18474 22480 32954 22536
rect 33010 22480 33015 22536
rect 18413 22478 33015 22480
rect 18413 22475 18479 22478
rect 32949 22475 33015 22478
rect 8170 22336 8486 22337
rect 8170 22272 8176 22336
rect 8240 22272 8256 22336
rect 8320 22272 8336 22336
rect 8400 22272 8416 22336
rect 8480 22272 8486 22336
rect 8170 22271 8486 22272
rect 22618 22336 22934 22337
rect 22618 22272 22624 22336
rect 22688 22272 22704 22336
rect 22768 22272 22784 22336
rect 22848 22272 22864 22336
rect 22928 22272 22934 22336
rect 22618 22271 22934 22272
rect 37066 22336 37382 22337
rect 37066 22272 37072 22336
rect 37136 22272 37152 22336
rect 37216 22272 37232 22336
rect 37296 22272 37312 22336
rect 37376 22272 37382 22336
rect 37066 22271 37382 22272
rect 51514 22336 51830 22337
rect 51514 22272 51520 22336
rect 51584 22272 51600 22336
rect 51664 22272 51680 22336
rect 51744 22272 51760 22336
rect 51824 22272 51830 22336
rect 51514 22271 51830 22272
rect 23933 22130 23999 22133
rect 24485 22130 24551 22133
rect 23933 22128 24551 22130
rect 23933 22072 23938 22128
rect 23994 22072 24490 22128
rect 24546 22072 24551 22128
rect 23933 22070 24551 22072
rect 23933 22067 23999 22070
rect 24485 22067 24551 22070
rect 19333 21994 19399 21997
rect 22093 21994 22159 21997
rect 22737 21994 22803 21997
rect 19333 21992 22803 21994
rect 19333 21936 19338 21992
rect 19394 21936 22098 21992
rect 22154 21936 22742 21992
rect 22798 21936 22803 21992
rect 19333 21934 22803 21936
rect 19333 21931 19399 21934
rect 22093 21931 22159 21934
rect 22737 21931 22803 21934
rect 47577 21994 47643 21997
rect 56593 21994 56659 21997
rect 47577 21992 56659 21994
rect 47577 21936 47582 21992
rect 47638 21936 56598 21992
rect 56654 21936 56659 21992
rect 47577 21934 56659 21936
rect 47577 21931 47643 21934
rect 56593 21931 56659 21934
rect 18873 21858 18939 21861
rect 21817 21858 21883 21861
rect 18873 21856 21883 21858
rect 18873 21800 18878 21856
rect 18934 21800 21822 21856
rect 21878 21800 21883 21856
rect 18873 21798 21883 21800
rect 18873 21795 18939 21798
rect 21817 21795 21883 21798
rect 15394 21792 15710 21793
rect 15394 21728 15400 21792
rect 15464 21728 15480 21792
rect 15544 21728 15560 21792
rect 15624 21728 15640 21792
rect 15704 21728 15710 21792
rect 15394 21727 15710 21728
rect 29842 21792 30158 21793
rect 29842 21728 29848 21792
rect 29912 21728 29928 21792
rect 29992 21728 30008 21792
rect 30072 21728 30088 21792
rect 30152 21728 30158 21792
rect 29842 21727 30158 21728
rect 44290 21792 44606 21793
rect 44290 21728 44296 21792
rect 44360 21728 44376 21792
rect 44440 21728 44456 21792
rect 44520 21728 44536 21792
rect 44600 21728 44606 21792
rect 44290 21727 44606 21728
rect 19425 21722 19491 21725
rect 25037 21722 25103 21725
rect 26141 21722 26207 21725
rect 19425 21720 26207 21722
rect 19425 21664 19430 21720
rect 19486 21664 25042 21720
rect 25098 21664 26146 21720
rect 26202 21664 26207 21720
rect 19425 21662 26207 21664
rect 19425 21659 19491 21662
rect 25037 21659 25103 21662
rect 26141 21659 26207 21662
rect 24485 21586 24551 21589
rect 27061 21586 27127 21589
rect 24485 21584 27127 21586
rect 24485 21528 24490 21584
rect 24546 21528 27066 21584
rect 27122 21528 27127 21584
rect 24485 21526 27127 21528
rect 24485 21523 24551 21526
rect 27061 21523 27127 21526
rect 29361 21450 29427 21453
rect 38009 21450 38075 21453
rect 29361 21448 38075 21450
rect 29361 21392 29366 21448
rect 29422 21392 38014 21448
rect 38070 21392 38075 21448
rect 29361 21390 38075 21392
rect 29361 21387 29427 21390
rect 38009 21387 38075 21390
rect 8170 21248 8486 21249
rect 8170 21184 8176 21248
rect 8240 21184 8256 21248
rect 8320 21184 8336 21248
rect 8400 21184 8416 21248
rect 8480 21184 8486 21248
rect 8170 21183 8486 21184
rect 22618 21248 22934 21249
rect 22618 21184 22624 21248
rect 22688 21184 22704 21248
rect 22768 21184 22784 21248
rect 22848 21184 22864 21248
rect 22928 21184 22934 21248
rect 22618 21183 22934 21184
rect 37066 21248 37382 21249
rect 37066 21184 37072 21248
rect 37136 21184 37152 21248
rect 37216 21184 37232 21248
rect 37296 21184 37312 21248
rect 37376 21184 37382 21248
rect 37066 21183 37382 21184
rect 51514 21248 51830 21249
rect 51514 21184 51520 21248
rect 51584 21184 51600 21248
rect 51664 21184 51680 21248
rect 51744 21184 51760 21248
rect 51824 21184 51830 21248
rect 51514 21183 51830 21184
rect 21541 21042 21607 21045
rect 36721 21042 36787 21045
rect 21541 21040 36787 21042
rect 21541 20984 21546 21040
rect 21602 20984 36726 21040
rect 36782 20984 36787 21040
rect 21541 20982 36787 20984
rect 21541 20979 21607 20982
rect 36721 20979 36787 20982
rect 15394 20704 15710 20705
rect 15394 20640 15400 20704
rect 15464 20640 15480 20704
rect 15544 20640 15560 20704
rect 15624 20640 15640 20704
rect 15704 20640 15710 20704
rect 15394 20639 15710 20640
rect 29842 20704 30158 20705
rect 29842 20640 29848 20704
rect 29912 20640 29928 20704
rect 29992 20640 30008 20704
rect 30072 20640 30088 20704
rect 30152 20640 30158 20704
rect 29842 20639 30158 20640
rect 44290 20704 44606 20705
rect 44290 20640 44296 20704
rect 44360 20640 44376 20704
rect 44440 20640 44456 20704
rect 44520 20640 44536 20704
rect 44600 20640 44606 20704
rect 44290 20639 44606 20640
rect 24301 20634 24367 20637
rect 28257 20634 28323 20637
rect 24301 20632 28323 20634
rect 24301 20576 24306 20632
rect 24362 20576 28262 20632
rect 28318 20576 28323 20632
rect 24301 20574 28323 20576
rect 24301 20571 24367 20574
rect 28257 20571 28323 20574
rect 0 20498 800 20528
rect 2957 20498 3023 20501
rect 0 20496 3023 20498
rect 0 20440 2962 20496
rect 3018 20440 3023 20496
rect 0 20438 3023 20440
rect 0 20408 800 20438
rect 2957 20435 3023 20438
rect 8170 20160 8486 20161
rect 8170 20096 8176 20160
rect 8240 20096 8256 20160
rect 8320 20096 8336 20160
rect 8400 20096 8416 20160
rect 8480 20096 8486 20160
rect 8170 20095 8486 20096
rect 22618 20160 22934 20161
rect 22618 20096 22624 20160
rect 22688 20096 22704 20160
rect 22768 20096 22784 20160
rect 22848 20096 22864 20160
rect 22928 20096 22934 20160
rect 22618 20095 22934 20096
rect 37066 20160 37382 20161
rect 37066 20096 37072 20160
rect 37136 20096 37152 20160
rect 37216 20096 37232 20160
rect 37296 20096 37312 20160
rect 37376 20096 37382 20160
rect 37066 20095 37382 20096
rect 51514 20160 51830 20161
rect 51514 20096 51520 20160
rect 51584 20096 51600 20160
rect 51664 20096 51680 20160
rect 51744 20096 51760 20160
rect 51824 20096 51830 20160
rect 51514 20095 51830 20096
rect 15837 20090 15903 20093
rect 22185 20090 22251 20093
rect 15837 20088 22251 20090
rect 15837 20032 15842 20088
rect 15898 20032 22190 20088
rect 22246 20032 22251 20088
rect 15837 20030 22251 20032
rect 15837 20027 15903 20030
rect 22185 20027 22251 20030
rect 18413 19954 18479 19957
rect 41781 19954 41847 19957
rect 18413 19952 41847 19954
rect 18413 19896 18418 19952
rect 18474 19896 41786 19952
rect 41842 19896 41847 19952
rect 18413 19894 41847 19896
rect 18413 19891 18479 19894
rect 41781 19891 41847 19894
rect 16573 19818 16639 19821
rect 19609 19818 19675 19821
rect 16573 19816 19675 19818
rect 16573 19760 16578 19816
rect 16634 19760 19614 19816
rect 19670 19760 19675 19816
rect 16573 19758 19675 19760
rect 16573 19755 16639 19758
rect 19609 19755 19675 19758
rect 19885 19818 19951 19821
rect 39205 19818 39271 19821
rect 19885 19816 39271 19818
rect 19885 19760 19890 19816
rect 19946 19760 39210 19816
rect 39266 19760 39271 19816
rect 19885 19758 39271 19760
rect 19885 19755 19951 19758
rect 39205 19755 39271 19758
rect 16481 19682 16547 19685
rect 27245 19682 27311 19685
rect 16481 19680 27311 19682
rect 16481 19624 16486 19680
rect 16542 19624 27250 19680
rect 27306 19624 27311 19680
rect 16481 19622 27311 19624
rect 16481 19619 16547 19622
rect 27245 19619 27311 19622
rect 15394 19616 15710 19617
rect 15394 19552 15400 19616
rect 15464 19552 15480 19616
rect 15544 19552 15560 19616
rect 15624 19552 15640 19616
rect 15704 19552 15710 19616
rect 15394 19551 15710 19552
rect 29842 19616 30158 19617
rect 29842 19552 29848 19616
rect 29912 19552 29928 19616
rect 29992 19552 30008 19616
rect 30072 19552 30088 19616
rect 30152 19552 30158 19616
rect 29842 19551 30158 19552
rect 44290 19616 44606 19617
rect 44290 19552 44296 19616
rect 44360 19552 44376 19616
rect 44440 19552 44456 19616
rect 44520 19552 44536 19616
rect 44600 19552 44606 19616
rect 44290 19551 44606 19552
rect 8170 19072 8486 19073
rect 8170 19008 8176 19072
rect 8240 19008 8256 19072
rect 8320 19008 8336 19072
rect 8400 19008 8416 19072
rect 8480 19008 8486 19072
rect 8170 19007 8486 19008
rect 22618 19072 22934 19073
rect 22618 19008 22624 19072
rect 22688 19008 22704 19072
rect 22768 19008 22784 19072
rect 22848 19008 22864 19072
rect 22928 19008 22934 19072
rect 22618 19007 22934 19008
rect 37066 19072 37382 19073
rect 37066 19008 37072 19072
rect 37136 19008 37152 19072
rect 37216 19008 37232 19072
rect 37296 19008 37312 19072
rect 37376 19008 37382 19072
rect 37066 19007 37382 19008
rect 51514 19072 51830 19073
rect 51514 19008 51520 19072
rect 51584 19008 51600 19072
rect 51664 19008 51680 19072
rect 51744 19008 51760 19072
rect 51824 19008 51830 19072
rect 51514 19007 51830 19008
rect 19241 18730 19307 18733
rect 33593 18730 33659 18733
rect 19241 18728 33659 18730
rect 19241 18672 19246 18728
rect 19302 18672 33598 18728
rect 33654 18672 33659 18728
rect 19241 18670 33659 18672
rect 19241 18667 19307 18670
rect 33593 18667 33659 18670
rect 15394 18528 15710 18529
rect 15394 18464 15400 18528
rect 15464 18464 15480 18528
rect 15544 18464 15560 18528
rect 15624 18464 15640 18528
rect 15704 18464 15710 18528
rect 15394 18463 15710 18464
rect 29842 18528 30158 18529
rect 29842 18464 29848 18528
rect 29912 18464 29928 18528
rect 29992 18464 30008 18528
rect 30072 18464 30088 18528
rect 30152 18464 30158 18528
rect 29842 18463 30158 18464
rect 44290 18528 44606 18529
rect 44290 18464 44296 18528
rect 44360 18464 44376 18528
rect 44440 18464 44456 18528
rect 44520 18464 44536 18528
rect 44600 18464 44606 18528
rect 44290 18463 44606 18464
rect 16021 18458 16087 18461
rect 18689 18458 18755 18461
rect 16021 18456 18755 18458
rect 16021 18400 16026 18456
rect 16082 18400 18694 18456
rect 18750 18400 18755 18456
rect 16021 18398 18755 18400
rect 16021 18395 16087 18398
rect 18689 18395 18755 18398
rect 3969 18322 4035 18325
rect 22185 18322 22251 18325
rect 22369 18322 22435 18325
rect 3969 18320 22435 18322
rect 3969 18264 3974 18320
rect 4030 18264 22190 18320
rect 22246 18264 22374 18320
rect 22430 18264 22435 18320
rect 3969 18262 22435 18264
rect 3969 18259 4035 18262
rect 22185 18259 22251 18262
rect 22369 18259 22435 18262
rect 27337 18322 27403 18325
rect 46841 18322 46907 18325
rect 27337 18320 46907 18322
rect 27337 18264 27342 18320
rect 27398 18264 46846 18320
rect 46902 18264 46907 18320
rect 27337 18262 46907 18264
rect 27337 18259 27403 18262
rect 46841 18259 46907 18262
rect 4061 18186 4127 18189
rect 14549 18186 14615 18189
rect 4061 18184 14615 18186
rect 4061 18128 4066 18184
rect 4122 18128 14554 18184
rect 14610 18128 14615 18184
rect 4061 18126 14615 18128
rect 4061 18123 4127 18126
rect 14549 18123 14615 18126
rect 38837 18186 38903 18189
rect 43345 18186 43411 18189
rect 38837 18184 43411 18186
rect 38837 18128 38842 18184
rect 38898 18128 43350 18184
rect 43406 18128 43411 18184
rect 38837 18126 43411 18128
rect 38837 18123 38903 18126
rect 43345 18123 43411 18126
rect 17769 18050 17835 18053
rect 22369 18050 22435 18053
rect 17769 18048 22435 18050
rect 17769 17992 17774 18048
rect 17830 17992 22374 18048
rect 22430 17992 22435 18048
rect 17769 17990 22435 17992
rect 17769 17987 17835 17990
rect 22369 17987 22435 17990
rect 8170 17984 8486 17985
rect 8170 17920 8176 17984
rect 8240 17920 8256 17984
rect 8320 17920 8336 17984
rect 8400 17920 8416 17984
rect 8480 17920 8486 17984
rect 8170 17919 8486 17920
rect 22618 17984 22934 17985
rect 22618 17920 22624 17984
rect 22688 17920 22704 17984
rect 22768 17920 22784 17984
rect 22848 17920 22864 17984
rect 22928 17920 22934 17984
rect 22618 17919 22934 17920
rect 37066 17984 37382 17985
rect 37066 17920 37072 17984
rect 37136 17920 37152 17984
rect 37216 17920 37232 17984
rect 37296 17920 37312 17984
rect 37376 17920 37382 17984
rect 37066 17919 37382 17920
rect 51514 17984 51830 17985
rect 51514 17920 51520 17984
rect 51584 17920 51600 17984
rect 51664 17920 51680 17984
rect 51744 17920 51760 17984
rect 51824 17920 51830 17984
rect 51514 17919 51830 17920
rect 51901 17914 51967 17917
rect 53833 17914 53899 17917
rect 51901 17912 53899 17914
rect 51901 17856 51906 17912
rect 51962 17856 53838 17912
rect 53894 17856 53899 17912
rect 51901 17854 53899 17856
rect 51901 17851 52010 17854
rect 53833 17851 53899 17854
rect 9305 17778 9371 17781
rect 48313 17778 48379 17781
rect 51950 17778 52010 17851
rect 9305 17776 52010 17778
rect 9305 17720 9310 17776
rect 9366 17720 48318 17776
rect 48374 17720 52010 17776
rect 9305 17718 52010 17720
rect 57789 17778 57855 17781
rect 59200 17778 60000 17808
rect 57789 17776 60000 17778
rect 57789 17720 57794 17776
rect 57850 17720 60000 17776
rect 57789 17718 60000 17720
rect 9305 17715 9371 17718
rect 48313 17715 48379 17718
rect 57789 17715 57855 17718
rect 59200 17688 60000 17718
rect 15101 17642 15167 17645
rect 31201 17642 31267 17645
rect 15101 17640 31267 17642
rect 15101 17584 15106 17640
rect 15162 17584 31206 17640
rect 31262 17584 31267 17640
rect 15101 17582 31267 17584
rect 15101 17579 15167 17582
rect 31201 17579 31267 17582
rect 32029 17642 32095 17645
rect 38101 17642 38167 17645
rect 32029 17640 38167 17642
rect 32029 17584 32034 17640
rect 32090 17584 38106 17640
rect 38162 17584 38167 17640
rect 32029 17582 38167 17584
rect 32029 17579 32095 17582
rect 38101 17579 38167 17582
rect 15394 17440 15710 17441
rect 15394 17376 15400 17440
rect 15464 17376 15480 17440
rect 15544 17376 15560 17440
rect 15624 17376 15640 17440
rect 15704 17376 15710 17440
rect 15394 17375 15710 17376
rect 29842 17440 30158 17441
rect 29842 17376 29848 17440
rect 29912 17376 29928 17440
rect 29992 17376 30008 17440
rect 30072 17376 30088 17440
rect 30152 17376 30158 17440
rect 29842 17375 30158 17376
rect 44290 17440 44606 17441
rect 44290 17376 44296 17440
rect 44360 17376 44376 17440
rect 44440 17376 44456 17440
rect 44520 17376 44536 17440
rect 44600 17376 44606 17440
rect 44290 17375 44606 17376
rect 21817 17370 21883 17373
rect 28349 17370 28415 17373
rect 21817 17368 28415 17370
rect 21817 17312 21822 17368
rect 21878 17312 28354 17368
rect 28410 17312 28415 17368
rect 21817 17310 28415 17312
rect 21817 17307 21883 17310
rect 28349 17307 28415 17310
rect 14917 17234 14983 17237
rect 23289 17234 23355 17237
rect 14917 17232 23355 17234
rect 14917 17176 14922 17232
rect 14978 17176 23294 17232
rect 23350 17176 23355 17232
rect 14917 17174 23355 17176
rect 14917 17171 14983 17174
rect 23289 17171 23355 17174
rect 38653 17234 38719 17237
rect 45185 17234 45251 17237
rect 38653 17232 45251 17234
rect 38653 17176 38658 17232
rect 38714 17176 45190 17232
rect 45246 17176 45251 17232
rect 38653 17174 45251 17176
rect 38653 17171 38719 17174
rect 45185 17171 45251 17174
rect 12065 17098 12131 17101
rect 21173 17098 21239 17101
rect 12065 17096 21239 17098
rect 12065 17040 12070 17096
rect 12126 17040 21178 17096
rect 21234 17040 21239 17096
rect 12065 17038 21239 17040
rect 12065 17035 12131 17038
rect 21173 17035 21239 17038
rect 26785 17098 26851 17101
rect 57237 17098 57303 17101
rect 26785 17096 57303 17098
rect 26785 17040 26790 17096
rect 26846 17040 57242 17096
rect 57298 17040 57303 17096
rect 26785 17038 57303 17040
rect 26785 17035 26851 17038
rect 57237 17035 57303 17038
rect 8170 16896 8486 16897
rect 8170 16832 8176 16896
rect 8240 16832 8256 16896
rect 8320 16832 8336 16896
rect 8400 16832 8416 16896
rect 8480 16832 8486 16896
rect 8170 16831 8486 16832
rect 22618 16896 22934 16897
rect 22618 16832 22624 16896
rect 22688 16832 22704 16896
rect 22768 16832 22784 16896
rect 22848 16832 22864 16896
rect 22928 16832 22934 16896
rect 22618 16831 22934 16832
rect 37066 16896 37382 16897
rect 37066 16832 37072 16896
rect 37136 16832 37152 16896
rect 37216 16832 37232 16896
rect 37296 16832 37312 16896
rect 37376 16832 37382 16896
rect 37066 16831 37382 16832
rect 51514 16896 51830 16897
rect 51514 16832 51520 16896
rect 51584 16832 51600 16896
rect 51664 16832 51680 16896
rect 51744 16832 51760 16896
rect 51824 16832 51830 16896
rect 51514 16831 51830 16832
rect 14089 16690 14155 16693
rect 34053 16690 34119 16693
rect 14089 16688 34119 16690
rect 14089 16632 14094 16688
rect 14150 16632 34058 16688
rect 34114 16632 34119 16688
rect 14089 16630 34119 16632
rect 14089 16627 14155 16630
rect 34053 16627 34119 16630
rect 6269 16554 6335 16557
rect 17217 16554 17283 16557
rect 6269 16552 17283 16554
rect 6269 16496 6274 16552
rect 6330 16496 17222 16552
rect 17278 16496 17283 16552
rect 6269 16494 17283 16496
rect 6269 16491 6335 16494
rect 17217 16491 17283 16494
rect 15394 16352 15710 16353
rect 15394 16288 15400 16352
rect 15464 16288 15480 16352
rect 15544 16288 15560 16352
rect 15624 16288 15640 16352
rect 15704 16288 15710 16352
rect 15394 16287 15710 16288
rect 29842 16352 30158 16353
rect 29842 16288 29848 16352
rect 29912 16288 29928 16352
rect 29992 16288 30008 16352
rect 30072 16288 30088 16352
rect 30152 16288 30158 16352
rect 29842 16287 30158 16288
rect 44290 16352 44606 16353
rect 44290 16288 44296 16352
rect 44360 16288 44376 16352
rect 44440 16288 44456 16352
rect 44520 16288 44536 16352
rect 44600 16288 44606 16352
rect 44290 16287 44606 16288
rect 4613 16282 4679 16285
rect 9121 16282 9187 16285
rect 4613 16280 9187 16282
rect 4613 16224 4618 16280
rect 4674 16224 9126 16280
rect 9182 16224 9187 16280
rect 4613 16222 9187 16224
rect 4613 16219 4679 16222
rect 9121 16219 9187 16222
rect 19701 16282 19767 16285
rect 29545 16282 29611 16285
rect 19701 16280 29611 16282
rect 19701 16224 19706 16280
rect 19762 16224 29550 16280
rect 29606 16224 29611 16280
rect 19701 16222 29611 16224
rect 19701 16219 19767 16222
rect 29545 16219 29611 16222
rect 4889 16146 4955 16149
rect 32121 16146 32187 16149
rect 4889 16144 32187 16146
rect 4889 16088 4894 16144
rect 4950 16088 32126 16144
rect 32182 16088 32187 16144
rect 4889 16086 32187 16088
rect 4889 16083 4955 16086
rect 32121 16083 32187 16086
rect 6453 16010 6519 16013
rect 18689 16010 18755 16013
rect 6453 16008 18755 16010
rect 6453 15952 6458 16008
rect 6514 15952 18694 16008
rect 18750 15952 18755 16008
rect 6453 15950 18755 15952
rect 6453 15947 6519 15950
rect 18689 15947 18755 15950
rect 20069 16010 20135 16013
rect 29637 16010 29703 16013
rect 20069 16008 29703 16010
rect 20069 15952 20074 16008
rect 20130 15952 29642 16008
rect 29698 15952 29703 16008
rect 20069 15950 29703 15952
rect 20069 15947 20135 15950
rect 29637 15947 29703 15950
rect 51165 16010 51231 16013
rect 57053 16010 57119 16013
rect 51165 16008 57119 16010
rect 51165 15952 51170 16008
rect 51226 15952 57058 16008
rect 57114 15952 57119 16008
rect 51165 15950 57119 15952
rect 51165 15947 51231 15950
rect 57053 15947 57119 15950
rect 8170 15808 8486 15809
rect 8170 15744 8176 15808
rect 8240 15744 8256 15808
rect 8320 15744 8336 15808
rect 8400 15744 8416 15808
rect 8480 15744 8486 15808
rect 8170 15743 8486 15744
rect 22618 15808 22934 15809
rect 22618 15744 22624 15808
rect 22688 15744 22704 15808
rect 22768 15744 22784 15808
rect 22848 15744 22864 15808
rect 22928 15744 22934 15808
rect 22618 15743 22934 15744
rect 37066 15808 37382 15809
rect 37066 15744 37072 15808
rect 37136 15744 37152 15808
rect 37216 15744 37232 15808
rect 37296 15744 37312 15808
rect 37376 15744 37382 15808
rect 37066 15743 37382 15744
rect 51514 15808 51830 15809
rect 51514 15744 51520 15808
rect 51584 15744 51600 15808
rect 51664 15744 51680 15808
rect 51744 15744 51760 15808
rect 51824 15744 51830 15808
rect 51514 15743 51830 15744
rect 38561 15738 38627 15741
rect 39113 15738 39179 15741
rect 41597 15738 41663 15741
rect 38561 15736 41663 15738
rect 38561 15680 38566 15736
rect 38622 15680 39118 15736
rect 39174 15680 41602 15736
rect 41658 15680 41663 15736
rect 38561 15678 41663 15680
rect 38561 15675 38627 15678
rect 39113 15675 39179 15678
rect 41597 15675 41663 15678
rect 8293 15602 8359 15605
rect 20897 15602 20963 15605
rect 8293 15600 20963 15602
rect 8293 15544 8298 15600
rect 8354 15544 20902 15600
rect 20958 15544 20963 15600
rect 8293 15542 20963 15544
rect 8293 15539 8359 15542
rect 20897 15539 20963 15542
rect 5717 15466 5783 15469
rect 28993 15466 29059 15469
rect 5717 15464 29059 15466
rect 5717 15408 5722 15464
rect 5778 15408 28998 15464
rect 29054 15408 29059 15464
rect 5717 15406 29059 15408
rect 5717 15403 5783 15406
rect 28993 15403 29059 15406
rect 50613 15466 50679 15469
rect 50981 15466 51047 15469
rect 52821 15466 52887 15469
rect 50613 15464 52887 15466
rect 50613 15408 50618 15464
rect 50674 15408 50986 15464
rect 51042 15408 52826 15464
rect 52882 15408 52887 15464
rect 50613 15406 52887 15408
rect 50613 15403 50679 15406
rect 50981 15403 51047 15406
rect 52821 15403 52887 15406
rect 15394 15264 15710 15265
rect 15394 15200 15400 15264
rect 15464 15200 15480 15264
rect 15544 15200 15560 15264
rect 15624 15200 15640 15264
rect 15704 15200 15710 15264
rect 15394 15199 15710 15200
rect 29842 15264 30158 15265
rect 29842 15200 29848 15264
rect 29912 15200 29928 15264
rect 29992 15200 30008 15264
rect 30072 15200 30088 15264
rect 30152 15200 30158 15264
rect 29842 15199 30158 15200
rect 44290 15264 44606 15265
rect 44290 15200 44296 15264
rect 44360 15200 44376 15264
rect 44440 15200 44456 15264
rect 44520 15200 44536 15264
rect 44600 15200 44606 15264
rect 44290 15199 44606 15200
rect 0 15058 800 15088
rect 21633 15058 21699 15061
rect 28809 15058 28875 15061
rect 0 14998 2790 15058
rect 0 14968 800 14998
rect 2730 13834 2790 14998
rect 21633 15056 28875 15058
rect 21633 15000 21638 15056
rect 21694 15000 28814 15056
rect 28870 15000 28875 15056
rect 21633 14998 28875 15000
rect 21633 14995 21699 14998
rect 28809 14995 28875 14998
rect 5441 14922 5507 14925
rect 17493 14922 17559 14925
rect 5441 14920 17559 14922
rect 5441 14864 5446 14920
rect 5502 14864 17498 14920
rect 17554 14864 17559 14920
rect 5441 14862 17559 14864
rect 5441 14859 5507 14862
rect 17493 14859 17559 14862
rect 8170 14720 8486 14721
rect 8170 14656 8176 14720
rect 8240 14656 8256 14720
rect 8320 14656 8336 14720
rect 8400 14656 8416 14720
rect 8480 14656 8486 14720
rect 8170 14655 8486 14656
rect 22618 14720 22934 14721
rect 22618 14656 22624 14720
rect 22688 14656 22704 14720
rect 22768 14656 22784 14720
rect 22848 14656 22864 14720
rect 22928 14656 22934 14720
rect 22618 14655 22934 14656
rect 37066 14720 37382 14721
rect 37066 14656 37072 14720
rect 37136 14656 37152 14720
rect 37216 14656 37232 14720
rect 37296 14656 37312 14720
rect 37376 14656 37382 14720
rect 37066 14655 37382 14656
rect 51514 14720 51830 14721
rect 51514 14656 51520 14720
rect 51584 14656 51600 14720
rect 51664 14656 51680 14720
rect 51744 14656 51760 14720
rect 51824 14656 51830 14720
rect 51514 14655 51830 14656
rect 8293 14514 8359 14517
rect 18965 14514 19031 14517
rect 8293 14512 19031 14514
rect 8293 14456 8298 14512
rect 8354 14456 18970 14512
rect 19026 14456 19031 14512
rect 8293 14454 19031 14456
rect 8293 14451 8359 14454
rect 18965 14451 19031 14454
rect 3785 14378 3851 14381
rect 16573 14378 16639 14381
rect 22001 14378 22067 14381
rect 3785 14376 22067 14378
rect 3785 14320 3790 14376
rect 3846 14320 16578 14376
rect 16634 14320 22006 14376
rect 22062 14320 22067 14376
rect 3785 14318 22067 14320
rect 3785 14315 3851 14318
rect 16573 14315 16639 14318
rect 22001 14315 22067 14318
rect 15394 14176 15710 14177
rect 15394 14112 15400 14176
rect 15464 14112 15480 14176
rect 15544 14112 15560 14176
rect 15624 14112 15640 14176
rect 15704 14112 15710 14176
rect 15394 14111 15710 14112
rect 29842 14176 30158 14177
rect 29842 14112 29848 14176
rect 29912 14112 29928 14176
rect 29992 14112 30008 14176
rect 30072 14112 30088 14176
rect 30152 14112 30158 14176
rect 29842 14111 30158 14112
rect 44290 14176 44606 14177
rect 44290 14112 44296 14176
rect 44360 14112 44376 14176
rect 44440 14112 44456 14176
rect 44520 14112 44536 14176
rect 44600 14112 44606 14176
rect 44290 14111 44606 14112
rect 20989 14106 21055 14109
rect 27613 14106 27679 14109
rect 20989 14104 27679 14106
rect 20989 14048 20994 14104
rect 21050 14048 27618 14104
rect 27674 14048 27679 14104
rect 20989 14046 27679 14048
rect 20989 14043 21055 14046
rect 27613 14043 27679 14046
rect 8753 13970 8819 13973
rect 30925 13970 30991 13973
rect 8753 13968 30991 13970
rect 8753 13912 8758 13968
rect 8814 13912 30930 13968
rect 30986 13912 30991 13968
rect 8753 13910 30991 13912
rect 8753 13907 8819 13910
rect 30925 13907 30991 13910
rect 18137 13834 18203 13837
rect 2730 13832 18203 13834
rect 2730 13776 18142 13832
rect 18198 13776 18203 13832
rect 2730 13774 18203 13776
rect 18137 13771 18203 13774
rect 8170 13632 8486 13633
rect 8170 13568 8176 13632
rect 8240 13568 8256 13632
rect 8320 13568 8336 13632
rect 8400 13568 8416 13632
rect 8480 13568 8486 13632
rect 8170 13567 8486 13568
rect 22618 13632 22934 13633
rect 22618 13568 22624 13632
rect 22688 13568 22704 13632
rect 22768 13568 22784 13632
rect 22848 13568 22864 13632
rect 22928 13568 22934 13632
rect 22618 13567 22934 13568
rect 37066 13632 37382 13633
rect 37066 13568 37072 13632
rect 37136 13568 37152 13632
rect 37216 13568 37232 13632
rect 37296 13568 37312 13632
rect 37376 13568 37382 13632
rect 37066 13567 37382 13568
rect 51514 13632 51830 13633
rect 51514 13568 51520 13632
rect 51584 13568 51600 13632
rect 51664 13568 51680 13632
rect 51744 13568 51760 13632
rect 51824 13568 51830 13632
rect 51514 13567 51830 13568
rect 6453 13290 6519 13293
rect 17309 13290 17375 13293
rect 6453 13288 17375 13290
rect 6453 13232 6458 13288
rect 6514 13232 17314 13288
rect 17370 13232 17375 13288
rect 6453 13230 17375 13232
rect 6453 13227 6519 13230
rect 17309 13227 17375 13230
rect 15394 13088 15710 13089
rect 15394 13024 15400 13088
rect 15464 13024 15480 13088
rect 15544 13024 15560 13088
rect 15624 13024 15640 13088
rect 15704 13024 15710 13088
rect 15394 13023 15710 13024
rect 29842 13088 30158 13089
rect 29842 13024 29848 13088
rect 29912 13024 29928 13088
rect 29992 13024 30008 13088
rect 30072 13024 30088 13088
rect 30152 13024 30158 13088
rect 29842 13023 30158 13024
rect 44290 13088 44606 13089
rect 44290 13024 44296 13088
rect 44360 13024 44376 13088
rect 44440 13024 44456 13088
rect 44520 13024 44536 13088
rect 44600 13024 44606 13088
rect 44290 13023 44606 13024
rect 58065 13018 58131 13021
rect 59200 13018 60000 13048
rect 58065 13016 60000 13018
rect 58065 12960 58070 13016
rect 58126 12960 60000 13016
rect 58065 12958 60000 12960
rect 58065 12955 58131 12958
rect 59200 12928 60000 12958
rect 12617 12882 12683 12885
rect 29821 12882 29887 12885
rect 12617 12880 29887 12882
rect 12617 12824 12622 12880
rect 12678 12824 29826 12880
rect 29882 12824 29887 12880
rect 12617 12822 29887 12824
rect 12617 12819 12683 12822
rect 29821 12819 29887 12822
rect 8170 12544 8486 12545
rect 8170 12480 8176 12544
rect 8240 12480 8256 12544
rect 8320 12480 8336 12544
rect 8400 12480 8416 12544
rect 8480 12480 8486 12544
rect 8170 12479 8486 12480
rect 22618 12544 22934 12545
rect 22618 12480 22624 12544
rect 22688 12480 22704 12544
rect 22768 12480 22784 12544
rect 22848 12480 22864 12544
rect 22928 12480 22934 12544
rect 22618 12479 22934 12480
rect 37066 12544 37382 12545
rect 37066 12480 37072 12544
rect 37136 12480 37152 12544
rect 37216 12480 37232 12544
rect 37296 12480 37312 12544
rect 37376 12480 37382 12544
rect 37066 12479 37382 12480
rect 51514 12544 51830 12545
rect 51514 12480 51520 12544
rect 51584 12480 51600 12544
rect 51664 12480 51680 12544
rect 51744 12480 51760 12544
rect 51824 12480 51830 12544
rect 51514 12479 51830 12480
rect 5809 12338 5875 12341
rect 22277 12338 22343 12341
rect 26877 12338 26943 12341
rect 5809 12336 22110 12338
rect 5809 12280 5814 12336
rect 5870 12280 22110 12336
rect 5809 12278 22110 12280
rect 5809 12275 5875 12278
rect 16389 12202 16455 12205
rect 18321 12202 18387 12205
rect 16389 12200 18387 12202
rect 16389 12144 16394 12200
rect 16450 12144 18326 12200
rect 18382 12144 18387 12200
rect 16389 12142 18387 12144
rect 22050 12202 22110 12278
rect 22277 12336 26943 12338
rect 22277 12280 22282 12336
rect 22338 12280 26882 12336
rect 26938 12280 26943 12336
rect 22277 12278 26943 12280
rect 22277 12275 22343 12278
rect 26877 12275 26943 12278
rect 26141 12202 26207 12205
rect 22050 12200 26207 12202
rect 22050 12144 26146 12200
rect 26202 12144 26207 12200
rect 22050 12142 26207 12144
rect 16389 12139 16455 12142
rect 18321 12139 18387 12142
rect 26141 12139 26207 12142
rect 15394 12000 15710 12001
rect 15394 11936 15400 12000
rect 15464 11936 15480 12000
rect 15544 11936 15560 12000
rect 15624 11936 15640 12000
rect 15704 11936 15710 12000
rect 15394 11935 15710 11936
rect 29842 12000 30158 12001
rect 29842 11936 29848 12000
rect 29912 11936 29928 12000
rect 29992 11936 30008 12000
rect 30072 11936 30088 12000
rect 30152 11936 30158 12000
rect 29842 11935 30158 11936
rect 44290 12000 44606 12001
rect 44290 11936 44296 12000
rect 44360 11936 44376 12000
rect 44440 11936 44456 12000
rect 44520 11936 44536 12000
rect 44600 11936 44606 12000
rect 44290 11935 44606 11936
rect 13537 11794 13603 11797
rect 23473 11794 23539 11797
rect 13537 11792 23539 11794
rect 13537 11736 13542 11792
rect 13598 11736 23478 11792
rect 23534 11736 23539 11792
rect 13537 11734 23539 11736
rect 13537 11731 13603 11734
rect 23473 11731 23539 11734
rect 19425 11658 19491 11661
rect 30373 11658 30439 11661
rect 30925 11658 30991 11661
rect 19425 11656 30991 11658
rect 19425 11600 19430 11656
rect 19486 11600 30378 11656
rect 30434 11600 30930 11656
rect 30986 11600 30991 11656
rect 19425 11598 30991 11600
rect 19425 11595 19491 11598
rect 30373 11595 30439 11598
rect 30925 11595 30991 11598
rect 8170 11456 8486 11457
rect 8170 11392 8176 11456
rect 8240 11392 8256 11456
rect 8320 11392 8336 11456
rect 8400 11392 8416 11456
rect 8480 11392 8486 11456
rect 8170 11391 8486 11392
rect 22618 11456 22934 11457
rect 22618 11392 22624 11456
rect 22688 11392 22704 11456
rect 22768 11392 22784 11456
rect 22848 11392 22864 11456
rect 22928 11392 22934 11456
rect 22618 11391 22934 11392
rect 37066 11456 37382 11457
rect 37066 11392 37072 11456
rect 37136 11392 37152 11456
rect 37216 11392 37232 11456
rect 37296 11392 37312 11456
rect 37376 11392 37382 11456
rect 37066 11391 37382 11392
rect 51514 11456 51830 11457
rect 51514 11392 51520 11456
rect 51584 11392 51600 11456
rect 51664 11392 51680 11456
rect 51744 11392 51760 11456
rect 51824 11392 51830 11456
rect 51514 11391 51830 11392
rect 38101 11114 38167 11117
rect 57605 11114 57671 11117
rect 38101 11112 57671 11114
rect 38101 11056 38106 11112
rect 38162 11056 57610 11112
rect 57666 11056 57671 11112
rect 38101 11054 57671 11056
rect 38101 11051 38167 11054
rect 57605 11051 57671 11054
rect 15394 10912 15710 10913
rect 15394 10848 15400 10912
rect 15464 10848 15480 10912
rect 15544 10848 15560 10912
rect 15624 10848 15640 10912
rect 15704 10848 15710 10912
rect 15394 10847 15710 10848
rect 29842 10912 30158 10913
rect 29842 10848 29848 10912
rect 29912 10848 29928 10912
rect 29992 10848 30008 10912
rect 30072 10848 30088 10912
rect 30152 10848 30158 10912
rect 29842 10847 30158 10848
rect 44290 10912 44606 10913
rect 44290 10848 44296 10912
rect 44360 10848 44376 10912
rect 44440 10848 44456 10912
rect 44520 10848 44536 10912
rect 44600 10848 44606 10912
rect 44290 10847 44606 10848
rect 37733 10706 37799 10709
rect 38469 10706 38535 10709
rect 37733 10704 38535 10706
rect 37733 10648 37738 10704
rect 37794 10648 38474 10704
rect 38530 10648 38535 10704
rect 37733 10646 38535 10648
rect 37733 10643 37799 10646
rect 38469 10643 38535 10646
rect 8170 10368 8486 10369
rect 0 10298 800 10328
rect 8170 10304 8176 10368
rect 8240 10304 8256 10368
rect 8320 10304 8336 10368
rect 8400 10304 8416 10368
rect 8480 10304 8486 10368
rect 8170 10303 8486 10304
rect 22618 10368 22934 10369
rect 22618 10304 22624 10368
rect 22688 10304 22704 10368
rect 22768 10304 22784 10368
rect 22848 10304 22864 10368
rect 22928 10304 22934 10368
rect 22618 10303 22934 10304
rect 37066 10368 37382 10369
rect 37066 10304 37072 10368
rect 37136 10304 37152 10368
rect 37216 10304 37232 10368
rect 37296 10304 37312 10368
rect 37376 10304 37382 10368
rect 37066 10303 37382 10304
rect 51514 10368 51830 10369
rect 51514 10304 51520 10368
rect 51584 10304 51600 10368
rect 51664 10304 51680 10368
rect 51744 10304 51760 10368
rect 51824 10304 51830 10368
rect 51514 10303 51830 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10208 800 10238
rect 1577 10235 1643 10238
rect 30465 10162 30531 10165
rect 36905 10162 36971 10165
rect 30465 10160 36971 10162
rect 30465 10104 30470 10160
rect 30526 10104 36910 10160
rect 36966 10104 36971 10160
rect 30465 10102 36971 10104
rect 30465 10099 30531 10102
rect 36905 10099 36971 10102
rect 21909 10026 21975 10029
rect 38653 10026 38719 10029
rect 21909 10024 38719 10026
rect 21909 9968 21914 10024
rect 21970 9968 38658 10024
rect 38714 9968 38719 10024
rect 21909 9966 38719 9968
rect 21909 9963 21975 9966
rect 38653 9963 38719 9966
rect 30281 9890 30347 9893
rect 31661 9890 31727 9893
rect 30281 9888 31727 9890
rect 30281 9832 30286 9888
rect 30342 9832 31666 9888
rect 31722 9832 31727 9888
rect 30281 9830 31727 9832
rect 30281 9827 30347 9830
rect 31661 9827 31727 9830
rect 15394 9824 15710 9825
rect 15394 9760 15400 9824
rect 15464 9760 15480 9824
rect 15544 9760 15560 9824
rect 15624 9760 15640 9824
rect 15704 9760 15710 9824
rect 15394 9759 15710 9760
rect 29842 9824 30158 9825
rect 29842 9760 29848 9824
rect 29912 9760 29928 9824
rect 29992 9760 30008 9824
rect 30072 9760 30088 9824
rect 30152 9760 30158 9824
rect 29842 9759 30158 9760
rect 44290 9824 44606 9825
rect 44290 9760 44296 9824
rect 44360 9760 44376 9824
rect 44440 9760 44456 9824
rect 44520 9760 44536 9824
rect 44600 9760 44606 9824
rect 44290 9759 44606 9760
rect 18413 9618 18479 9621
rect 55397 9618 55463 9621
rect 18413 9616 55463 9618
rect 18413 9560 18418 9616
rect 18474 9560 55402 9616
rect 55458 9560 55463 9616
rect 18413 9558 55463 9560
rect 18413 9555 18479 9558
rect 55397 9555 55463 9558
rect 8170 9280 8486 9281
rect 8170 9216 8176 9280
rect 8240 9216 8256 9280
rect 8320 9216 8336 9280
rect 8400 9216 8416 9280
rect 8480 9216 8486 9280
rect 8170 9215 8486 9216
rect 22618 9280 22934 9281
rect 22618 9216 22624 9280
rect 22688 9216 22704 9280
rect 22768 9216 22784 9280
rect 22848 9216 22864 9280
rect 22928 9216 22934 9280
rect 22618 9215 22934 9216
rect 37066 9280 37382 9281
rect 37066 9216 37072 9280
rect 37136 9216 37152 9280
rect 37216 9216 37232 9280
rect 37296 9216 37312 9280
rect 37376 9216 37382 9280
rect 37066 9215 37382 9216
rect 51514 9280 51830 9281
rect 51514 9216 51520 9280
rect 51584 9216 51600 9280
rect 51664 9216 51680 9280
rect 51744 9216 51760 9280
rect 51824 9216 51830 9280
rect 51514 9215 51830 9216
rect 29729 9074 29795 9077
rect 32765 9074 32831 9077
rect 29729 9072 32831 9074
rect 29729 9016 29734 9072
rect 29790 9016 32770 9072
rect 32826 9016 32831 9072
rect 29729 9014 32831 9016
rect 29729 9011 29795 9014
rect 32765 9011 32831 9014
rect 21173 8938 21239 8941
rect 55581 8938 55647 8941
rect 21173 8936 55647 8938
rect 21173 8880 21178 8936
rect 21234 8880 55586 8936
rect 55642 8880 55647 8936
rect 21173 8878 55647 8880
rect 21173 8875 21239 8878
rect 55581 8875 55647 8878
rect 15394 8736 15710 8737
rect 15394 8672 15400 8736
rect 15464 8672 15480 8736
rect 15544 8672 15560 8736
rect 15624 8672 15640 8736
rect 15704 8672 15710 8736
rect 15394 8671 15710 8672
rect 29842 8736 30158 8737
rect 29842 8672 29848 8736
rect 29912 8672 29928 8736
rect 29992 8672 30008 8736
rect 30072 8672 30088 8736
rect 30152 8672 30158 8736
rect 29842 8671 30158 8672
rect 44290 8736 44606 8737
rect 44290 8672 44296 8736
rect 44360 8672 44376 8736
rect 44440 8672 44456 8736
rect 44520 8672 44536 8736
rect 44600 8672 44606 8736
rect 44290 8671 44606 8672
rect 38653 8666 38719 8669
rect 40861 8666 40927 8669
rect 38653 8664 40927 8666
rect 38653 8608 38658 8664
rect 38714 8608 40866 8664
rect 40922 8608 40927 8664
rect 38653 8606 40927 8608
rect 38653 8603 38719 8606
rect 40861 8603 40927 8606
rect 30925 8530 30991 8533
rect 39757 8530 39823 8533
rect 30925 8528 39823 8530
rect 30925 8472 30930 8528
rect 30986 8472 39762 8528
rect 39818 8472 39823 8528
rect 30925 8470 39823 8472
rect 30925 8467 30991 8470
rect 39757 8467 39823 8470
rect 39849 8394 39915 8397
rect 44817 8394 44883 8397
rect 39849 8392 44883 8394
rect 39849 8336 39854 8392
rect 39910 8336 44822 8392
rect 44878 8336 44883 8392
rect 39849 8334 44883 8336
rect 39849 8331 39915 8334
rect 44817 8331 44883 8334
rect 39665 8258 39731 8261
rect 43069 8258 43135 8261
rect 46381 8258 46447 8261
rect 39665 8256 46447 8258
rect 39665 8200 39670 8256
rect 39726 8200 43074 8256
rect 43130 8200 46386 8256
rect 46442 8200 46447 8256
rect 39665 8198 46447 8200
rect 39665 8195 39731 8198
rect 43069 8195 43135 8198
rect 46381 8195 46447 8198
rect 8170 8192 8486 8193
rect 8170 8128 8176 8192
rect 8240 8128 8256 8192
rect 8320 8128 8336 8192
rect 8400 8128 8416 8192
rect 8480 8128 8486 8192
rect 8170 8127 8486 8128
rect 22618 8192 22934 8193
rect 22618 8128 22624 8192
rect 22688 8128 22704 8192
rect 22768 8128 22784 8192
rect 22848 8128 22864 8192
rect 22928 8128 22934 8192
rect 22618 8127 22934 8128
rect 37066 8192 37382 8193
rect 37066 8128 37072 8192
rect 37136 8128 37152 8192
rect 37216 8128 37232 8192
rect 37296 8128 37312 8192
rect 37376 8128 37382 8192
rect 37066 8127 37382 8128
rect 51514 8192 51830 8193
rect 51514 8128 51520 8192
rect 51584 8128 51600 8192
rect 51664 8128 51680 8192
rect 51744 8128 51760 8192
rect 51824 8128 51830 8192
rect 51514 8127 51830 8128
rect 31109 8122 31175 8125
rect 31753 8122 31819 8125
rect 31109 8120 31819 8122
rect 31109 8064 31114 8120
rect 31170 8064 31758 8120
rect 31814 8064 31819 8120
rect 31109 8062 31819 8064
rect 31109 8059 31175 8062
rect 31753 8059 31819 8062
rect 31661 7986 31727 7989
rect 39021 7986 39087 7989
rect 31661 7984 39087 7986
rect 31661 7928 31666 7984
rect 31722 7928 39026 7984
rect 39082 7928 39087 7984
rect 31661 7926 39087 7928
rect 31661 7923 31727 7926
rect 39021 7923 39087 7926
rect 27797 7850 27863 7853
rect 33685 7850 33751 7853
rect 27797 7848 33751 7850
rect 27797 7792 27802 7848
rect 27858 7792 33690 7848
rect 33746 7792 33751 7848
rect 27797 7790 33751 7792
rect 27797 7787 27863 7790
rect 33685 7787 33751 7790
rect 15394 7648 15710 7649
rect 15394 7584 15400 7648
rect 15464 7584 15480 7648
rect 15544 7584 15560 7648
rect 15624 7584 15640 7648
rect 15704 7584 15710 7648
rect 15394 7583 15710 7584
rect 29842 7648 30158 7649
rect 29842 7584 29848 7648
rect 29912 7584 29928 7648
rect 29992 7584 30008 7648
rect 30072 7584 30088 7648
rect 30152 7584 30158 7648
rect 29842 7583 30158 7584
rect 44290 7648 44606 7649
rect 44290 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44536 7648
rect 44600 7584 44606 7648
rect 44290 7583 44606 7584
rect 58065 7578 58131 7581
rect 59200 7578 60000 7608
rect 58065 7576 60000 7578
rect 58065 7520 58070 7576
rect 58126 7520 60000 7576
rect 58065 7518 60000 7520
rect 58065 7515 58131 7518
rect 59200 7488 60000 7518
rect 28257 7442 28323 7445
rect 33041 7442 33107 7445
rect 28257 7440 33107 7442
rect 28257 7384 28262 7440
rect 28318 7384 33046 7440
rect 33102 7384 33107 7440
rect 28257 7382 33107 7384
rect 28257 7379 28323 7382
rect 33041 7379 33107 7382
rect 8170 7104 8486 7105
rect 8170 7040 8176 7104
rect 8240 7040 8256 7104
rect 8320 7040 8336 7104
rect 8400 7040 8416 7104
rect 8480 7040 8486 7104
rect 8170 7039 8486 7040
rect 22618 7104 22934 7105
rect 22618 7040 22624 7104
rect 22688 7040 22704 7104
rect 22768 7040 22784 7104
rect 22848 7040 22864 7104
rect 22928 7040 22934 7104
rect 22618 7039 22934 7040
rect 37066 7104 37382 7105
rect 37066 7040 37072 7104
rect 37136 7040 37152 7104
rect 37216 7040 37232 7104
rect 37296 7040 37312 7104
rect 37376 7040 37382 7104
rect 37066 7039 37382 7040
rect 51514 7104 51830 7105
rect 51514 7040 51520 7104
rect 51584 7040 51600 7104
rect 51664 7040 51680 7104
rect 51744 7040 51760 7104
rect 51824 7040 51830 7104
rect 51514 7039 51830 7040
rect 28809 7034 28875 7037
rect 30557 7034 30623 7037
rect 31109 7034 31175 7037
rect 31569 7034 31635 7037
rect 28809 7032 31635 7034
rect 28809 6976 28814 7032
rect 28870 6976 30562 7032
rect 30618 6976 31114 7032
rect 31170 6976 31574 7032
rect 31630 6976 31635 7032
rect 28809 6974 31635 6976
rect 28809 6971 28875 6974
rect 30557 6971 30623 6974
rect 31109 6971 31175 6974
rect 31569 6971 31635 6974
rect 31569 6898 31635 6901
rect 38285 6898 38351 6901
rect 31569 6896 38351 6898
rect 31569 6840 31574 6896
rect 31630 6840 38290 6896
rect 38346 6840 38351 6896
rect 31569 6838 38351 6840
rect 31569 6835 31635 6838
rect 38285 6835 38351 6838
rect 15394 6560 15710 6561
rect 15394 6496 15400 6560
rect 15464 6496 15480 6560
rect 15544 6496 15560 6560
rect 15624 6496 15640 6560
rect 15704 6496 15710 6560
rect 15394 6495 15710 6496
rect 29842 6560 30158 6561
rect 29842 6496 29848 6560
rect 29912 6496 29928 6560
rect 29992 6496 30008 6560
rect 30072 6496 30088 6560
rect 30152 6496 30158 6560
rect 29842 6495 30158 6496
rect 44290 6560 44606 6561
rect 44290 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44536 6560
rect 44600 6496 44606 6560
rect 44290 6495 44606 6496
rect 8170 6016 8486 6017
rect 8170 5952 8176 6016
rect 8240 5952 8256 6016
rect 8320 5952 8336 6016
rect 8400 5952 8416 6016
rect 8480 5952 8486 6016
rect 8170 5951 8486 5952
rect 22618 6016 22934 6017
rect 22618 5952 22624 6016
rect 22688 5952 22704 6016
rect 22768 5952 22784 6016
rect 22848 5952 22864 6016
rect 22928 5952 22934 6016
rect 22618 5951 22934 5952
rect 37066 6016 37382 6017
rect 37066 5952 37072 6016
rect 37136 5952 37152 6016
rect 37216 5952 37232 6016
rect 37296 5952 37312 6016
rect 37376 5952 37382 6016
rect 37066 5951 37382 5952
rect 51514 6016 51830 6017
rect 51514 5952 51520 6016
rect 51584 5952 51600 6016
rect 51664 5952 51680 6016
rect 51744 5952 51760 6016
rect 51824 5952 51830 6016
rect 51514 5951 51830 5952
rect 15394 5472 15710 5473
rect 15394 5408 15400 5472
rect 15464 5408 15480 5472
rect 15544 5408 15560 5472
rect 15624 5408 15640 5472
rect 15704 5408 15710 5472
rect 15394 5407 15710 5408
rect 29842 5472 30158 5473
rect 29842 5408 29848 5472
rect 29912 5408 29928 5472
rect 29992 5408 30008 5472
rect 30072 5408 30088 5472
rect 30152 5408 30158 5472
rect 29842 5407 30158 5408
rect 44290 5472 44606 5473
rect 44290 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44536 5472
rect 44600 5408 44606 5472
rect 44290 5407 44606 5408
rect 8170 4928 8486 4929
rect 0 4858 800 4888
rect 8170 4864 8176 4928
rect 8240 4864 8256 4928
rect 8320 4864 8336 4928
rect 8400 4864 8416 4928
rect 8480 4864 8486 4928
rect 8170 4863 8486 4864
rect 22618 4928 22934 4929
rect 22618 4864 22624 4928
rect 22688 4864 22704 4928
rect 22768 4864 22784 4928
rect 22848 4864 22864 4928
rect 22928 4864 22934 4928
rect 22618 4863 22934 4864
rect 37066 4928 37382 4929
rect 37066 4864 37072 4928
rect 37136 4864 37152 4928
rect 37216 4864 37232 4928
rect 37296 4864 37312 4928
rect 37376 4864 37382 4928
rect 37066 4863 37382 4864
rect 51514 4928 51830 4929
rect 51514 4864 51520 4928
rect 51584 4864 51600 4928
rect 51664 4864 51680 4928
rect 51744 4864 51760 4928
rect 51824 4864 51830 4928
rect 51514 4863 51830 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 24853 4586 24919 4589
rect 42057 4586 42123 4589
rect 24853 4584 42123 4586
rect 24853 4528 24858 4584
rect 24914 4528 42062 4584
rect 42118 4528 42123 4584
rect 24853 4526 42123 4528
rect 24853 4523 24919 4526
rect 42057 4523 42123 4526
rect 15394 4384 15710 4385
rect 15394 4320 15400 4384
rect 15464 4320 15480 4384
rect 15544 4320 15560 4384
rect 15624 4320 15640 4384
rect 15704 4320 15710 4384
rect 15394 4319 15710 4320
rect 29842 4384 30158 4385
rect 29842 4320 29848 4384
rect 29912 4320 29928 4384
rect 29992 4320 30008 4384
rect 30072 4320 30088 4384
rect 30152 4320 30158 4384
rect 29842 4319 30158 4320
rect 44290 4384 44606 4385
rect 44290 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44536 4384
rect 44600 4320 44606 4384
rect 44290 4319 44606 4320
rect 8170 3840 8486 3841
rect 8170 3776 8176 3840
rect 8240 3776 8256 3840
rect 8320 3776 8336 3840
rect 8400 3776 8416 3840
rect 8480 3776 8486 3840
rect 8170 3775 8486 3776
rect 22618 3840 22934 3841
rect 22618 3776 22624 3840
rect 22688 3776 22704 3840
rect 22768 3776 22784 3840
rect 22848 3776 22864 3840
rect 22928 3776 22934 3840
rect 22618 3775 22934 3776
rect 37066 3840 37382 3841
rect 37066 3776 37072 3840
rect 37136 3776 37152 3840
rect 37216 3776 37232 3840
rect 37296 3776 37312 3840
rect 37376 3776 37382 3840
rect 37066 3775 37382 3776
rect 51514 3840 51830 3841
rect 51514 3776 51520 3840
rect 51584 3776 51600 3840
rect 51664 3776 51680 3840
rect 51744 3776 51760 3840
rect 51824 3776 51830 3840
rect 51514 3775 51830 3776
rect 15394 3296 15710 3297
rect 15394 3232 15400 3296
rect 15464 3232 15480 3296
rect 15544 3232 15560 3296
rect 15624 3232 15640 3296
rect 15704 3232 15710 3296
rect 15394 3231 15710 3232
rect 29842 3296 30158 3297
rect 29842 3232 29848 3296
rect 29912 3232 29928 3296
rect 29992 3232 30008 3296
rect 30072 3232 30088 3296
rect 30152 3232 30158 3296
rect 29842 3231 30158 3232
rect 44290 3296 44606 3297
rect 44290 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44536 3296
rect 44600 3232 44606 3296
rect 44290 3231 44606 3232
rect 58065 2818 58131 2821
rect 59200 2818 60000 2848
rect 58065 2816 60000 2818
rect 58065 2760 58070 2816
rect 58126 2760 60000 2816
rect 58065 2758 60000 2760
rect 58065 2755 58131 2758
rect 8170 2752 8486 2753
rect 8170 2688 8176 2752
rect 8240 2688 8256 2752
rect 8320 2688 8336 2752
rect 8400 2688 8416 2752
rect 8480 2688 8486 2752
rect 8170 2687 8486 2688
rect 22618 2752 22934 2753
rect 22618 2688 22624 2752
rect 22688 2688 22704 2752
rect 22768 2688 22784 2752
rect 22848 2688 22864 2752
rect 22928 2688 22934 2752
rect 22618 2687 22934 2688
rect 37066 2752 37382 2753
rect 37066 2688 37072 2752
rect 37136 2688 37152 2752
rect 37216 2688 37232 2752
rect 37296 2688 37312 2752
rect 37376 2688 37382 2752
rect 37066 2687 37382 2688
rect 51514 2752 51830 2753
rect 51514 2688 51520 2752
rect 51584 2688 51600 2752
rect 51664 2688 51680 2752
rect 51744 2688 51760 2752
rect 51824 2688 51830 2752
rect 59200 2728 60000 2758
rect 51514 2687 51830 2688
rect 15394 2208 15710 2209
rect 15394 2144 15400 2208
rect 15464 2144 15480 2208
rect 15544 2144 15560 2208
rect 15624 2144 15640 2208
rect 15704 2144 15710 2208
rect 15394 2143 15710 2144
rect 29842 2208 30158 2209
rect 29842 2144 29848 2208
rect 29912 2144 29928 2208
rect 29992 2144 30008 2208
rect 30072 2144 30088 2208
rect 30152 2144 30158 2208
rect 29842 2143 30158 2144
rect 44290 2208 44606 2209
rect 44290 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44536 2208
rect 44600 2144 44606 2208
rect 44290 2143 44606 2144
<< via3 >>
rect 15400 33756 15464 33760
rect 15400 33700 15404 33756
rect 15404 33700 15460 33756
rect 15460 33700 15464 33756
rect 15400 33696 15464 33700
rect 15480 33756 15544 33760
rect 15480 33700 15484 33756
rect 15484 33700 15540 33756
rect 15540 33700 15544 33756
rect 15480 33696 15544 33700
rect 15560 33756 15624 33760
rect 15560 33700 15564 33756
rect 15564 33700 15620 33756
rect 15620 33700 15624 33756
rect 15560 33696 15624 33700
rect 15640 33756 15704 33760
rect 15640 33700 15644 33756
rect 15644 33700 15700 33756
rect 15700 33700 15704 33756
rect 15640 33696 15704 33700
rect 29848 33756 29912 33760
rect 29848 33700 29852 33756
rect 29852 33700 29908 33756
rect 29908 33700 29912 33756
rect 29848 33696 29912 33700
rect 29928 33756 29992 33760
rect 29928 33700 29932 33756
rect 29932 33700 29988 33756
rect 29988 33700 29992 33756
rect 29928 33696 29992 33700
rect 30008 33756 30072 33760
rect 30008 33700 30012 33756
rect 30012 33700 30068 33756
rect 30068 33700 30072 33756
rect 30008 33696 30072 33700
rect 30088 33756 30152 33760
rect 30088 33700 30092 33756
rect 30092 33700 30148 33756
rect 30148 33700 30152 33756
rect 30088 33696 30152 33700
rect 44296 33756 44360 33760
rect 44296 33700 44300 33756
rect 44300 33700 44356 33756
rect 44356 33700 44360 33756
rect 44296 33696 44360 33700
rect 44376 33756 44440 33760
rect 44376 33700 44380 33756
rect 44380 33700 44436 33756
rect 44436 33700 44440 33756
rect 44376 33696 44440 33700
rect 44456 33756 44520 33760
rect 44456 33700 44460 33756
rect 44460 33700 44516 33756
rect 44516 33700 44520 33756
rect 44456 33696 44520 33700
rect 44536 33756 44600 33760
rect 44536 33700 44540 33756
rect 44540 33700 44596 33756
rect 44596 33700 44600 33756
rect 44536 33696 44600 33700
rect 8176 33212 8240 33216
rect 8176 33156 8180 33212
rect 8180 33156 8236 33212
rect 8236 33156 8240 33212
rect 8176 33152 8240 33156
rect 8256 33212 8320 33216
rect 8256 33156 8260 33212
rect 8260 33156 8316 33212
rect 8316 33156 8320 33212
rect 8256 33152 8320 33156
rect 8336 33212 8400 33216
rect 8336 33156 8340 33212
rect 8340 33156 8396 33212
rect 8396 33156 8400 33212
rect 8336 33152 8400 33156
rect 8416 33212 8480 33216
rect 8416 33156 8420 33212
rect 8420 33156 8476 33212
rect 8476 33156 8480 33212
rect 8416 33152 8480 33156
rect 22624 33212 22688 33216
rect 22624 33156 22628 33212
rect 22628 33156 22684 33212
rect 22684 33156 22688 33212
rect 22624 33152 22688 33156
rect 22704 33212 22768 33216
rect 22704 33156 22708 33212
rect 22708 33156 22764 33212
rect 22764 33156 22768 33212
rect 22704 33152 22768 33156
rect 22784 33212 22848 33216
rect 22784 33156 22788 33212
rect 22788 33156 22844 33212
rect 22844 33156 22848 33212
rect 22784 33152 22848 33156
rect 22864 33212 22928 33216
rect 22864 33156 22868 33212
rect 22868 33156 22924 33212
rect 22924 33156 22928 33212
rect 22864 33152 22928 33156
rect 37072 33212 37136 33216
rect 37072 33156 37076 33212
rect 37076 33156 37132 33212
rect 37132 33156 37136 33212
rect 37072 33152 37136 33156
rect 37152 33212 37216 33216
rect 37152 33156 37156 33212
rect 37156 33156 37212 33212
rect 37212 33156 37216 33212
rect 37152 33152 37216 33156
rect 37232 33212 37296 33216
rect 37232 33156 37236 33212
rect 37236 33156 37292 33212
rect 37292 33156 37296 33212
rect 37232 33152 37296 33156
rect 37312 33212 37376 33216
rect 37312 33156 37316 33212
rect 37316 33156 37372 33212
rect 37372 33156 37376 33212
rect 37312 33152 37376 33156
rect 51520 33212 51584 33216
rect 51520 33156 51524 33212
rect 51524 33156 51580 33212
rect 51580 33156 51584 33212
rect 51520 33152 51584 33156
rect 51600 33212 51664 33216
rect 51600 33156 51604 33212
rect 51604 33156 51660 33212
rect 51660 33156 51664 33212
rect 51600 33152 51664 33156
rect 51680 33212 51744 33216
rect 51680 33156 51684 33212
rect 51684 33156 51740 33212
rect 51740 33156 51744 33212
rect 51680 33152 51744 33156
rect 51760 33212 51824 33216
rect 51760 33156 51764 33212
rect 51764 33156 51820 33212
rect 51820 33156 51824 33212
rect 51760 33152 51824 33156
rect 15400 32668 15464 32672
rect 15400 32612 15404 32668
rect 15404 32612 15460 32668
rect 15460 32612 15464 32668
rect 15400 32608 15464 32612
rect 15480 32668 15544 32672
rect 15480 32612 15484 32668
rect 15484 32612 15540 32668
rect 15540 32612 15544 32668
rect 15480 32608 15544 32612
rect 15560 32668 15624 32672
rect 15560 32612 15564 32668
rect 15564 32612 15620 32668
rect 15620 32612 15624 32668
rect 15560 32608 15624 32612
rect 15640 32668 15704 32672
rect 15640 32612 15644 32668
rect 15644 32612 15700 32668
rect 15700 32612 15704 32668
rect 15640 32608 15704 32612
rect 29848 32668 29912 32672
rect 29848 32612 29852 32668
rect 29852 32612 29908 32668
rect 29908 32612 29912 32668
rect 29848 32608 29912 32612
rect 29928 32668 29992 32672
rect 29928 32612 29932 32668
rect 29932 32612 29988 32668
rect 29988 32612 29992 32668
rect 29928 32608 29992 32612
rect 30008 32668 30072 32672
rect 30008 32612 30012 32668
rect 30012 32612 30068 32668
rect 30068 32612 30072 32668
rect 30008 32608 30072 32612
rect 30088 32668 30152 32672
rect 30088 32612 30092 32668
rect 30092 32612 30148 32668
rect 30148 32612 30152 32668
rect 30088 32608 30152 32612
rect 44296 32668 44360 32672
rect 44296 32612 44300 32668
rect 44300 32612 44356 32668
rect 44356 32612 44360 32668
rect 44296 32608 44360 32612
rect 44376 32668 44440 32672
rect 44376 32612 44380 32668
rect 44380 32612 44436 32668
rect 44436 32612 44440 32668
rect 44376 32608 44440 32612
rect 44456 32668 44520 32672
rect 44456 32612 44460 32668
rect 44460 32612 44516 32668
rect 44516 32612 44520 32668
rect 44456 32608 44520 32612
rect 44536 32668 44600 32672
rect 44536 32612 44540 32668
rect 44540 32612 44596 32668
rect 44596 32612 44600 32668
rect 44536 32608 44600 32612
rect 8176 32124 8240 32128
rect 8176 32068 8180 32124
rect 8180 32068 8236 32124
rect 8236 32068 8240 32124
rect 8176 32064 8240 32068
rect 8256 32124 8320 32128
rect 8256 32068 8260 32124
rect 8260 32068 8316 32124
rect 8316 32068 8320 32124
rect 8256 32064 8320 32068
rect 8336 32124 8400 32128
rect 8336 32068 8340 32124
rect 8340 32068 8396 32124
rect 8396 32068 8400 32124
rect 8336 32064 8400 32068
rect 8416 32124 8480 32128
rect 8416 32068 8420 32124
rect 8420 32068 8476 32124
rect 8476 32068 8480 32124
rect 8416 32064 8480 32068
rect 22624 32124 22688 32128
rect 22624 32068 22628 32124
rect 22628 32068 22684 32124
rect 22684 32068 22688 32124
rect 22624 32064 22688 32068
rect 22704 32124 22768 32128
rect 22704 32068 22708 32124
rect 22708 32068 22764 32124
rect 22764 32068 22768 32124
rect 22704 32064 22768 32068
rect 22784 32124 22848 32128
rect 22784 32068 22788 32124
rect 22788 32068 22844 32124
rect 22844 32068 22848 32124
rect 22784 32064 22848 32068
rect 22864 32124 22928 32128
rect 22864 32068 22868 32124
rect 22868 32068 22924 32124
rect 22924 32068 22928 32124
rect 22864 32064 22928 32068
rect 37072 32124 37136 32128
rect 37072 32068 37076 32124
rect 37076 32068 37132 32124
rect 37132 32068 37136 32124
rect 37072 32064 37136 32068
rect 37152 32124 37216 32128
rect 37152 32068 37156 32124
rect 37156 32068 37212 32124
rect 37212 32068 37216 32124
rect 37152 32064 37216 32068
rect 37232 32124 37296 32128
rect 37232 32068 37236 32124
rect 37236 32068 37292 32124
rect 37292 32068 37296 32124
rect 37232 32064 37296 32068
rect 37312 32124 37376 32128
rect 37312 32068 37316 32124
rect 37316 32068 37372 32124
rect 37372 32068 37376 32124
rect 37312 32064 37376 32068
rect 51520 32124 51584 32128
rect 51520 32068 51524 32124
rect 51524 32068 51580 32124
rect 51580 32068 51584 32124
rect 51520 32064 51584 32068
rect 51600 32124 51664 32128
rect 51600 32068 51604 32124
rect 51604 32068 51660 32124
rect 51660 32068 51664 32124
rect 51600 32064 51664 32068
rect 51680 32124 51744 32128
rect 51680 32068 51684 32124
rect 51684 32068 51740 32124
rect 51740 32068 51744 32124
rect 51680 32064 51744 32068
rect 51760 32124 51824 32128
rect 51760 32068 51764 32124
rect 51764 32068 51820 32124
rect 51820 32068 51824 32124
rect 51760 32064 51824 32068
rect 15400 31580 15464 31584
rect 15400 31524 15404 31580
rect 15404 31524 15460 31580
rect 15460 31524 15464 31580
rect 15400 31520 15464 31524
rect 15480 31580 15544 31584
rect 15480 31524 15484 31580
rect 15484 31524 15540 31580
rect 15540 31524 15544 31580
rect 15480 31520 15544 31524
rect 15560 31580 15624 31584
rect 15560 31524 15564 31580
rect 15564 31524 15620 31580
rect 15620 31524 15624 31580
rect 15560 31520 15624 31524
rect 15640 31580 15704 31584
rect 15640 31524 15644 31580
rect 15644 31524 15700 31580
rect 15700 31524 15704 31580
rect 15640 31520 15704 31524
rect 29848 31580 29912 31584
rect 29848 31524 29852 31580
rect 29852 31524 29908 31580
rect 29908 31524 29912 31580
rect 29848 31520 29912 31524
rect 29928 31580 29992 31584
rect 29928 31524 29932 31580
rect 29932 31524 29988 31580
rect 29988 31524 29992 31580
rect 29928 31520 29992 31524
rect 30008 31580 30072 31584
rect 30008 31524 30012 31580
rect 30012 31524 30068 31580
rect 30068 31524 30072 31580
rect 30008 31520 30072 31524
rect 30088 31580 30152 31584
rect 30088 31524 30092 31580
rect 30092 31524 30148 31580
rect 30148 31524 30152 31580
rect 30088 31520 30152 31524
rect 44296 31580 44360 31584
rect 44296 31524 44300 31580
rect 44300 31524 44356 31580
rect 44356 31524 44360 31580
rect 44296 31520 44360 31524
rect 44376 31580 44440 31584
rect 44376 31524 44380 31580
rect 44380 31524 44436 31580
rect 44436 31524 44440 31580
rect 44376 31520 44440 31524
rect 44456 31580 44520 31584
rect 44456 31524 44460 31580
rect 44460 31524 44516 31580
rect 44516 31524 44520 31580
rect 44456 31520 44520 31524
rect 44536 31580 44600 31584
rect 44536 31524 44540 31580
rect 44540 31524 44596 31580
rect 44596 31524 44600 31580
rect 44536 31520 44600 31524
rect 8176 31036 8240 31040
rect 8176 30980 8180 31036
rect 8180 30980 8236 31036
rect 8236 30980 8240 31036
rect 8176 30976 8240 30980
rect 8256 31036 8320 31040
rect 8256 30980 8260 31036
rect 8260 30980 8316 31036
rect 8316 30980 8320 31036
rect 8256 30976 8320 30980
rect 8336 31036 8400 31040
rect 8336 30980 8340 31036
rect 8340 30980 8396 31036
rect 8396 30980 8400 31036
rect 8336 30976 8400 30980
rect 8416 31036 8480 31040
rect 8416 30980 8420 31036
rect 8420 30980 8476 31036
rect 8476 30980 8480 31036
rect 8416 30976 8480 30980
rect 22624 31036 22688 31040
rect 22624 30980 22628 31036
rect 22628 30980 22684 31036
rect 22684 30980 22688 31036
rect 22624 30976 22688 30980
rect 22704 31036 22768 31040
rect 22704 30980 22708 31036
rect 22708 30980 22764 31036
rect 22764 30980 22768 31036
rect 22704 30976 22768 30980
rect 22784 31036 22848 31040
rect 22784 30980 22788 31036
rect 22788 30980 22844 31036
rect 22844 30980 22848 31036
rect 22784 30976 22848 30980
rect 22864 31036 22928 31040
rect 22864 30980 22868 31036
rect 22868 30980 22924 31036
rect 22924 30980 22928 31036
rect 22864 30976 22928 30980
rect 37072 31036 37136 31040
rect 37072 30980 37076 31036
rect 37076 30980 37132 31036
rect 37132 30980 37136 31036
rect 37072 30976 37136 30980
rect 37152 31036 37216 31040
rect 37152 30980 37156 31036
rect 37156 30980 37212 31036
rect 37212 30980 37216 31036
rect 37152 30976 37216 30980
rect 37232 31036 37296 31040
rect 37232 30980 37236 31036
rect 37236 30980 37292 31036
rect 37292 30980 37296 31036
rect 37232 30976 37296 30980
rect 37312 31036 37376 31040
rect 37312 30980 37316 31036
rect 37316 30980 37372 31036
rect 37372 30980 37376 31036
rect 37312 30976 37376 30980
rect 51520 31036 51584 31040
rect 51520 30980 51524 31036
rect 51524 30980 51580 31036
rect 51580 30980 51584 31036
rect 51520 30976 51584 30980
rect 51600 31036 51664 31040
rect 51600 30980 51604 31036
rect 51604 30980 51660 31036
rect 51660 30980 51664 31036
rect 51600 30976 51664 30980
rect 51680 31036 51744 31040
rect 51680 30980 51684 31036
rect 51684 30980 51740 31036
rect 51740 30980 51744 31036
rect 51680 30976 51744 30980
rect 51760 31036 51824 31040
rect 51760 30980 51764 31036
rect 51764 30980 51820 31036
rect 51820 30980 51824 31036
rect 51760 30976 51824 30980
rect 15400 30492 15464 30496
rect 15400 30436 15404 30492
rect 15404 30436 15460 30492
rect 15460 30436 15464 30492
rect 15400 30432 15464 30436
rect 15480 30492 15544 30496
rect 15480 30436 15484 30492
rect 15484 30436 15540 30492
rect 15540 30436 15544 30492
rect 15480 30432 15544 30436
rect 15560 30492 15624 30496
rect 15560 30436 15564 30492
rect 15564 30436 15620 30492
rect 15620 30436 15624 30492
rect 15560 30432 15624 30436
rect 15640 30492 15704 30496
rect 15640 30436 15644 30492
rect 15644 30436 15700 30492
rect 15700 30436 15704 30492
rect 15640 30432 15704 30436
rect 29848 30492 29912 30496
rect 29848 30436 29852 30492
rect 29852 30436 29908 30492
rect 29908 30436 29912 30492
rect 29848 30432 29912 30436
rect 29928 30492 29992 30496
rect 29928 30436 29932 30492
rect 29932 30436 29988 30492
rect 29988 30436 29992 30492
rect 29928 30432 29992 30436
rect 30008 30492 30072 30496
rect 30008 30436 30012 30492
rect 30012 30436 30068 30492
rect 30068 30436 30072 30492
rect 30008 30432 30072 30436
rect 30088 30492 30152 30496
rect 30088 30436 30092 30492
rect 30092 30436 30148 30492
rect 30148 30436 30152 30492
rect 30088 30432 30152 30436
rect 44296 30492 44360 30496
rect 44296 30436 44300 30492
rect 44300 30436 44356 30492
rect 44356 30436 44360 30492
rect 44296 30432 44360 30436
rect 44376 30492 44440 30496
rect 44376 30436 44380 30492
rect 44380 30436 44436 30492
rect 44436 30436 44440 30492
rect 44376 30432 44440 30436
rect 44456 30492 44520 30496
rect 44456 30436 44460 30492
rect 44460 30436 44516 30492
rect 44516 30436 44520 30492
rect 44456 30432 44520 30436
rect 44536 30492 44600 30496
rect 44536 30436 44540 30492
rect 44540 30436 44596 30492
rect 44596 30436 44600 30492
rect 44536 30432 44600 30436
rect 8176 29948 8240 29952
rect 8176 29892 8180 29948
rect 8180 29892 8236 29948
rect 8236 29892 8240 29948
rect 8176 29888 8240 29892
rect 8256 29948 8320 29952
rect 8256 29892 8260 29948
rect 8260 29892 8316 29948
rect 8316 29892 8320 29948
rect 8256 29888 8320 29892
rect 8336 29948 8400 29952
rect 8336 29892 8340 29948
rect 8340 29892 8396 29948
rect 8396 29892 8400 29948
rect 8336 29888 8400 29892
rect 8416 29948 8480 29952
rect 8416 29892 8420 29948
rect 8420 29892 8476 29948
rect 8476 29892 8480 29948
rect 8416 29888 8480 29892
rect 22624 29948 22688 29952
rect 22624 29892 22628 29948
rect 22628 29892 22684 29948
rect 22684 29892 22688 29948
rect 22624 29888 22688 29892
rect 22704 29948 22768 29952
rect 22704 29892 22708 29948
rect 22708 29892 22764 29948
rect 22764 29892 22768 29948
rect 22704 29888 22768 29892
rect 22784 29948 22848 29952
rect 22784 29892 22788 29948
rect 22788 29892 22844 29948
rect 22844 29892 22848 29948
rect 22784 29888 22848 29892
rect 22864 29948 22928 29952
rect 22864 29892 22868 29948
rect 22868 29892 22924 29948
rect 22924 29892 22928 29948
rect 22864 29888 22928 29892
rect 37072 29948 37136 29952
rect 37072 29892 37076 29948
rect 37076 29892 37132 29948
rect 37132 29892 37136 29948
rect 37072 29888 37136 29892
rect 37152 29948 37216 29952
rect 37152 29892 37156 29948
rect 37156 29892 37212 29948
rect 37212 29892 37216 29948
rect 37152 29888 37216 29892
rect 37232 29948 37296 29952
rect 37232 29892 37236 29948
rect 37236 29892 37292 29948
rect 37292 29892 37296 29948
rect 37232 29888 37296 29892
rect 37312 29948 37376 29952
rect 37312 29892 37316 29948
rect 37316 29892 37372 29948
rect 37372 29892 37376 29948
rect 37312 29888 37376 29892
rect 51520 29948 51584 29952
rect 51520 29892 51524 29948
rect 51524 29892 51580 29948
rect 51580 29892 51584 29948
rect 51520 29888 51584 29892
rect 51600 29948 51664 29952
rect 51600 29892 51604 29948
rect 51604 29892 51660 29948
rect 51660 29892 51664 29948
rect 51600 29888 51664 29892
rect 51680 29948 51744 29952
rect 51680 29892 51684 29948
rect 51684 29892 51740 29948
rect 51740 29892 51744 29948
rect 51680 29888 51744 29892
rect 51760 29948 51824 29952
rect 51760 29892 51764 29948
rect 51764 29892 51820 29948
rect 51820 29892 51824 29948
rect 51760 29888 51824 29892
rect 15400 29404 15464 29408
rect 15400 29348 15404 29404
rect 15404 29348 15460 29404
rect 15460 29348 15464 29404
rect 15400 29344 15464 29348
rect 15480 29404 15544 29408
rect 15480 29348 15484 29404
rect 15484 29348 15540 29404
rect 15540 29348 15544 29404
rect 15480 29344 15544 29348
rect 15560 29404 15624 29408
rect 15560 29348 15564 29404
rect 15564 29348 15620 29404
rect 15620 29348 15624 29404
rect 15560 29344 15624 29348
rect 15640 29404 15704 29408
rect 15640 29348 15644 29404
rect 15644 29348 15700 29404
rect 15700 29348 15704 29404
rect 15640 29344 15704 29348
rect 29848 29404 29912 29408
rect 29848 29348 29852 29404
rect 29852 29348 29908 29404
rect 29908 29348 29912 29404
rect 29848 29344 29912 29348
rect 29928 29404 29992 29408
rect 29928 29348 29932 29404
rect 29932 29348 29988 29404
rect 29988 29348 29992 29404
rect 29928 29344 29992 29348
rect 30008 29404 30072 29408
rect 30008 29348 30012 29404
rect 30012 29348 30068 29404
rect 30068 29348 30072 29404
rect 30008 29344 30072 29348
rect 30088 29404 30152 29408
rect 30088 29348 30092 29404
rect 30092 29348 30148 29404
rect 30148 29348 30152 29404
rect 30088 29344 30152 29348
rect 44296 29404 44360 29408
rect 44296 29348 44300 29404
rect 44300 29348 44356 29404
rect 44356 29348 44360 29404
rect 44296 29344 44360 29348
rect 44376 29404 44440 29408
rect 44376 29348 44380 29404
rect 44380 29348 44436 29404
rect 44436 29348 44440 29404
rect 44376 29344 44440 29348
rect 44456 29404 44520 29408
rect 44456 29348 44460 29404
rect 44460 29348 44516 29404
rect 44516 29348 44520 29404
rect 44456 29344 44520 29348
rect 44536 29404 44600 29408
rect 44536 29348 44540 29404
rect 44540 29348 44596 29404
rect 44596 29348 44600 29404
rect 44536 29344 44600 29348
rect 8176 28860 8240 28864
rect 8176 28804 8180 28860
rect 8180 28804 8236 28860
rect 8236 28804 8240 28860
rect 8176 28800 8240 28804
rect 8256 28860 8320 28864
rect 8256 28804 8260 28860
rect 8260 28804 8316 28860
rect 8316 28804 8320 28860
rect 8256 28800 8320 28804
rect 8336 28860 8400 28864
rect 8336 28804 8340 28860
rect 8340 28804 8396 28860
rect 8396 28804 8400 28860
rect 8336 28800 8400 28804
rect 8416 28860 8480 28864
rect 8416 28804 8420 28860
rect 8420 28804 8476 28860
rect 8476 28804 8480 28860
rect 8416 28800 8480 28804
rect 22624 28860 22688 28864
rect 22624 28804 22628 28860
rect 22628 28804 22684 28860
rect 22684 28804 22688 28860
rect 22624 28800 22688 28804
rect 22704 28860 22768 28864
rect 22704 28804 22708 28860
rect 22708 28804 22764 28860
rect 22764 28804 22768 28860
rect 22704 28800 22768 28804
rect 22784 28860 22848 28864
rect 22784 28804 22788 28860
rect 22788 28804 22844 28860
rect 22844 28804 22848 28860
rect 22784 28800 22848 28804
rect 22864 28860 22928 28864
rect 22864 28804 22868 28860
rect 22868 28804 22924 28860
rect 22924 28804 22928 28860
rect 22864 28800 22928 28804
rect 37072 28860 37136 28864
rect 37072 28804 37076 28860
rect 37076 28804 37132 28860
rect 37132 28804 37136 28860
rect 37072 28800 37136 28804
rect 37152 28860 37216 28864
rect 37152 28804 37156 28860
rect 37156 28804 37212 28860
rect 37212 28804 37216 28860
rect 37152 28800 37216 28804
rect 37232 28860 37296 28864
rect 37232 28804 37236 28860
rect 37236 28804 37292 28860
rect 37292 28804 37296 28860
rect 37232 28800 37296 28804
rect 37312 28860 37376 28864
rect 37312 28804 37316 28860
rect 37316 28804 37372 28860
rect 37372 28804 37376 28860
rect 37312 28800 37376 28804
rect 51520 28860 51584 28864
rect 51520 28804 51524 28860
rect 51524 28804 51580 28860
rect 51580 28804 51584 28860
rect 51520 28800 51584 28804
rect 51600 28860 51664 28864
rect 51600 28804 51604 28860
rect 51604 28804 51660 28860
rect 51660 28804 51664 28860
rect 51600 28800 51664 28804
rect 51680 28860 51744 28864
rect 51680 28804 51684 28860
rect 51684 28804 51740 28860
rect 51740 28804 51744 28860
rect 51680 28800 51744 28804
rect 51760 28860 51824 28864
rect 51760 28804 51764 28860
rect 51764 28804 51820 28860
rect 51820 28804 51824 28860
rect 51760 28800 51824 28804
rect 15400 28316 15464 28320
rect 15400 28260 15404 28316
rect 15404 28260 15460 28316
rect 15460 28260 15464 28316
rect 15400 28256 15464 28260
rect 15480 28316 15544 28320
rect 15480 28260 15484 28316
rect 15484 28260 15540 28316
rect 15540 28260 15544 28316
rect 15480 28256 15544 28260
rect 15560 28316 15624 28320
rect 15560 28260 15564 28316
rect 15564 28260 15620 28316
rect 15620 28260 15624 28316
rect 15560 28256 15624 28260
rect 15640 28316 15704 28320
rect 15640 28260 15644 28316
rect 15644 28260 15700 28316
rect 15700 28260 15704 28316
rect 15640 28256 15704 28260
rect 29848 28316 29912 28320
rect 29848 28260 29852 28316
rect 29852 28260 29908 28316
rect 29908 28260 29912 28316
rect 29848 28256 29912 28260
rect 29928 28316 29992 28320
rect 29928 28260 29932 28316
rect 29932 28260 29988 28316
rect 29988 28260 29992 28316
rect 29928 28256 29992 28260
rect 30008 28316 30072 28320
rect 30008 28260 30012 28316
rect 30012 28260 30068 28316
rect 30068 28260 30072 28316
rect 30008 28256 30072 28260
rect 30088 28316 30152 28320
rect 30088 28260 30092 28316
rect 30092 28260 30148 28316
rect 30148 28260 30152 28316
rect 30088 28256 30152 28260
rect 44296 28316 44360 28320
rect 44296 28260 44300 28316
rect 44300 28260 44356 28316
rect 44356 28260 44360 28316
rect 44296 28256 44360 28260
rect 44376 28316 44440 28320
rect 44376 28260 44380 28316
rect 44380 28260 44436 28316
rect 44436 28260 44440 28316
rect 44376 28256 44440 28260
rect 44456 28316 44520 28320
rect 44456 28260 44460 28316
rect 44460 28260 44516 28316
rect 44516 28260 44520 28316
rect 44456 28256 44520 28260
rect 44536 28316 44600 28320
rect 44536 28260 44540 28316
rect 44540 28260 44596 28316
rect 44596 28260 44600 28316
rect 44536 28256 44600 28260
rect 8176 27772 8240 27776
rect 8176 27716 8180 27772
rect 8180 27716 8236 27772
rect 8236 27716 8240 27772
rect 8176 27712 8240 27716
rect 8256 27772 8320 27776
rect 8256 27716 8260 27772
rect 8260 27716 8316 27772
rect 8316 27716 8320 27772
rect 8256 27712 8320 27716
rect 8336 27772 8400 27776
rect 8336 27716 8340 27772
rect 8340 27716 8396 27772
rect 8396 27716 8400 27772
rect 8336 27712 8400 27716
rect 8416 27772 8480 27776
rect 8416 27716 8420 27772
rect 8420 27716 8476 27772
rect 8476 27716 8480 27772
rect 8416 27712 8480 27716
rect 22624 27772 22688 27776
rect 22624 27716 22628 27772
rect 22628 27716 22684 27772
rect 22684 27716 22688 27772
rect 22624 27712 22688 27716
rect 22704 27772 22768 27776
rect 22704 27716 22708 27772
rect 22708 27716 22764 27772
rect 22764 27716 22768 27772
rect 22704 27712 22768 27716
rect 22784 27772 22848 27776
rect 22784 27716 22788 27772
rect 22788 27716 22844 27772
rect 22844 27716 22848 27772
rect 22784 27712 22848 27716
rect 22864 27772 22928 27776
rect 22864 27716 22868 27772
rect 22868 27716 22924 27772
rect 22924 27716 22928 27772
rect 22864 27712 22928 27716
rect 37072 27772 37136 27776
rect 37072 27716 37076 27772
rect 37076 27716 37132 27772
rect 37132 27716 37136 27772
rect 37072 27712 37136 27716
rect 37152 27772 37216 27776
rect 37152 27716 37156 27772
rect 37156 27716 37212 27772
rect 37212 27716 37216 27772
rect 37152 27712 37216 27716
rect 37232 27772 37296 27776
rect 37232 27716 37236 27772
rect 37236 27716 37292 27772
rect 37292 27716 37296 27772
rect 37232 27712 37296 27716
rect 37312 27772 37376 27776
rect 37312 27716 37316 27772
rect 37316 27716 37372 27772
rect 37372 27716 37376 27772
rect 37312 27712 37376 27716
rect 51520 27772 51584 27776
rect 51520 27716 51524 27772
rect 51524 27716 51580 27772
rect 51580 27716 51584 27772
rect 51520 27712 51584 27716
rect 51600 27772 51664 27776
rect 51600 27716 51604 27772
rect 51604 27716 51660 27772
rect 51660 27716 51664 27772
rect 51600 27712 51664 27716
rect 51680 27772 51744 27776
rect 51680 27716 51684 27772
rect 51684 27716 51740 27772
rect 51740 27716 51744 27772
rect 51680 27712 51744 27716
rect 51760 27772 51824 27776
rect 51760 27716 51764 27772
rect 51764 27716 51820 27772
rect 51820 27716 51824 27772
rect 51760 27712 51824 27716
rect 15400 27228 15464 27232
rect 15400 27172 15404 27228
rect 15404 27172 15460 27228
rect 15460 27172 15464 27228
rect 15400 27168 15464 27172
rect 15480 27228 15544 27232
rect 15480 27172 15484 27228
rect 15484 27172 15540 27228
rect 15540 27172 15544 27228
rect 15480 27168 15544 27172
rect 15560 27228 15624 27232
rect 15560 27172 15564 27228
rect 15564 27172 15620 27228
rect 15620 27172 15624 27228
rect 15560 27168 15624 27172
rect 15640 27228 15704 27232
rect 15640 27172 15644 27228
rect 15644 27172 15700 27228
rect 15700 27172 15704 27228
rect 15640 27168 15704 27172
rect 29848 27228 29912 27232
rect 29848 27172 29852 27228
rect 29852 27172 29908 27228
rect 29908 27172 29912 27228
rect 29848 27168 29912 27172
rect 29928 27228 29992 27232
rect 29928 27172 29932 27228
rect 29932 27172 29988 27228
rect 29988 27172 29992 27228
rect 29928 27168 29992 27172
rect 30008 27228 30072 27232
rect 30008 27172 30012 27228
rect 30012 27172 30068 27228
rect 30068 27172 30072 27228
rect 30008 27168 30072 27172
rect 30088 27228 30152 27232
rect 30088 27172 30092 27228
rect 30092 27172 30148 27228
rect 30148 27172 30152 27228
rect 30088 27168 30152 27172
rect 44296 27228 44360 27232
rect 44296 27172 44300 27228
rect 44300 27172 44356 27228
rect 44356 27172 44360 27228
rect 44296 27168 44360 27172
rect 44376 27228 44440 27232
rect 44376 27172 44380 27228
rect 44380 27172 44436 27228
rect 44436 27172 44440 27228
rect 44376 27168 44440 27172
rect 44456 27228 44520 27232
rect 44456 27172 44460 27228
rect 44460 27172 44516 27228
rect 44516 27172 44520 27228
rect 44456 27168 44520 27172
rect 44536 27228 44600 27232
rect 44536 27172 44540 27228
rect 44540 27172 44596 27228
rect 44596 27172 44600 27228
rect 44536 27168 44600 27172
rect 8176 26684 8240 26688
rect 8176 26628 8180 26684
rect 8180 26628 8236 26684
rect 8236 26628 8240 26684
rect 8176 26624 8240 26628
rect 8256 26684 8320 26688
rect 8256 26628 8260 26684
rect 8260 26628 8316 26684
rect 8316 26628 8320 26684
rect 8256 26624 8320 26628
rect 8336 26684 8400 26688
rect 8336 26628 8340 26684
rect 8340 26628 8396 26684
rect 8396 26628 8400 26684
rect 8336 26624 8400 26628
rect 8416 26684 8480 26688
rect 8416 26628 8420 26684
rect 8420 26628 8476 26684
rect 8476 26628 8480 26684
rect 8416 26624 8480 26628
rect 22624 26684 22688 26688
rect 22624 26628 22628 26684
rect 22628 26628 22684 26684
rect 22684 26628 22688 26684
rect 22624 26624 22688 26628
rect 22704 26684 22768 26688
rect 22704 26628 22708 26684
rect 22708 26628 22764 26684
rect 22764 26628 22768 26684
rect 22704 26624 22768 26628
rect 22784 26684 22848 26688
rect 22784 26628 22788 26684
rect 22788 26628 22844 26684
rect 22844 26628 22848 26684
rect 22784 26624 22848 26628
rect 22864 26684 22928 26688
rect 22864 26628 22868 26684
rect 22868 26628 22924 26684
rect 22924 26628 22928 26684
rect 22864 26624 22928 26628
rect 37072 26684 37136 26688
rect 37072 26628 37076 26684
rect 37076 26628 37132 26684
rect 37132 26628 37136 26684
rect 37072 26624 37136 26628
rect 37152 26684 37216 26688
rect 37152 26628 37156 26684
rect 37156 26628 37212 26684
rect 37212 26628 37216 26684
rect 37152 26624 37216 26628
rect 37232 26684 37296 26688
rect 37232 26628 37236 26684
rect 37236 26628 37292 26684
rect 37292 26628 37296 26684
rect 37232 26624 37296 26628
rect 37312 26684 37376 26688
rect 37312 26628 37316 26684
rect 37316 26628 37372 26684
rect 37372 26628 37376 26684
rect 37312 26624 37376 26628
rect 51520 26684 51584 26688
rect 51520 26628 51524 26684
rect 51524 26628 51580 26684
rect 51580 26628 51584 26684
rect 51520 26624 51584 26628
rect 51600 26684 51664 26688
rect 51600 26628 51604 26684
rect 51604 26628 51660 26684
rect 51660 26628 51664 26684
rect 51600 26624 51664 26628
rect 51680 26684 51744 26688
rect 51680 26628 51684 26684
rect 51684 26628 51740 26684
rect 51740 26628 51744 26684
rect 51680 26624 51744 26628
rect 51760 26684 51824 26688
rect 51760 26628 51764 26684
rect 51764 26628 51820 26684
rect 51820 26628 51824 26684
rect 51760 26624 51824 26628
rect 15400 26140 15464 26144
rect 15400 26084 15404 26140
rect 15404 26084 15460 26140
rect 15460 26084 15464 26140
rect 15400 26080 15464 26084
rect 15480 26140 15544 26144
rect 15480 26084 15484 26140
rect 15484 26084 15540 26140
rect 15540 26084 15544 26140
rect 15480 26080 15544 26084
rect 15560 26140 15624 26144
rect 15560 26084 15564 26140
rect 15564 26084 15620 26140
rect 15620 26084 15624 26140
rect 15560 26080 15624 26084
rect 15640 26140 15704 26144
rect 15640 26084 15644 26140
rect 15644 26084 15700 26140
rect 15700 26084 15704 26140
rect 15640 26080 15704 26084
rect 29848 26140 29912 26144
rect 29848 26084 29852 26140
rect 29852 26084 29908 26140
rect 29908 26084 29912 26140
rect 29848 26080 29912 26084
rect 29928 26140 29992 26144
rect 29928 26084 29932 26140
rect 29932 26084 29988 26140
rect 29988 26084 29992 26140
rect 29928 26080 29992 26084
rect 30008 26140 30072 26144
rect 30008 26084 30012 26140
rect 30012 26084 30068 26140
rect 30068 26084 30072 26140
rect 30008 26080 30072 26084
rect 30088 26140 30152 26144
rect 30088 26084 30092 26140
rect 30092 26084 30148 26140
rect 30148 26084 30152 26140
rect 30088 26080 30152 26084
rect 44296 26140 44360 26144
rect 44296 26084 44300 26140
rect 44300 26084 44356 26140
rect 44356 26084 44360 26140
rect 44296 26080 44360 26084
rect 44376 26140 44440 26144
rect 44376 26084 44380 26140
rect 44380 26084 44436 26140
rect 44436 26084 44440 26140
rect 44376 26080 44440 26084
rect 44456 26140 44520 26144
rect 44456 26084 44460 26140
rect 44460 26084 44516 26140
rect 44516 26084 44520 26140
rect 44456 26080 44520 26084
rect 44536 26140 44600 26144
rect 44536 26084 44540 26140
rect 44540 26084 44596 26140
rect 44596 26084 44600 26140
rect 44536 26080 44600 26084
rect 8176 25596 8240 25600
rect 8176 25540 8180 25596
rect 8180 25540 8236 25596
rect 8236 25540 8240 25596
rect 8176 25536 8240 25540
rect 8256 25596 8320 25600
rect 8256 25540 8260 25596
rect 8260 25540 8316 25596
rect 8316 25540 8320 25596
rect 8256 25536 8320 25540
rect 8336 25596 8400 25600
rect 8336 25540 8340 25596
rect 8340 25540 8396 25596
rect 8396 25540 8400 25596
rect 8336 25536 8400 25540
rect 8416 25596 8480 25600
rect 8416 25540 8420 25596
rect 8420 25540 8476 25596
rect 8476 25540 8480 25596
rect 8416 25536 8480 25540
rect 22624 25596 22688 25600
rect 22624 25540 22628 25596
rect 22628 25540 22684 25596
rect 22684 25540 22688 25596
rect 22624 25536 22688 25540
rect 22704 25596 22768 25600
rect 22704 25540 22708 25596
rect 22708 25540 22764 25596
rect 22764 25540 22768 25596
rect 22704 25536 22768 25540
rect 22784 25596 22848 25600
rect 22784 25540 22788 25596
rect 22788 25540 22844 25596
rect 22844 25540 22848 25596
rect 22784 25536 22848 25540
rect 22864 25596 22928 25600
rect 22864 25540 22868 25596
rect 22868 25540 22924 25596
rect 22924 25540 22928 25596
rect 22864 25536 22928 25540
rect 37072 25596 37136 25600
rect 37072 25540 37076 25596
rect 37076 25540 37132 25596
rect 37132 25540 37136 25596
rect 37072 25536 37136 25540
rect 37152 25596 37216 25600
rect 37152 25540 37156 25596
rect 37156 25540 37212 25596
rect 37212 25540 37216 25596
rect 37152 25536 37216 25540
rect 37232 25596 37296 25600
rect 37232 25540 37236 25596
rect 37236 25540 37292 25596
rect 37292 25540 37296 25596
rect 37232 25536 37296 25540
rect 37312 25596 37376 25600
rect 37312 25540 37316 25596
rect 37316 25540 37372 25596
rect 37372 25540 37376 25596
rect 37312 25536 37376 25540
rect 51520 25596 51584 25600
rect 51520 25540 51524 25596
rect 51524 25540 51580 25596
rect 51580 25540 51584 25596
rect 51520 25536 51584 25540
rect 51600 25596 51664 25600
rect 51600 25540 51604 25596
rect 51604 25540 51660 25596
rect 51660 25540 51664 25596
rect 51600 25536 51664 25540
rect 51680 25596 51744 25600
rect 51680 25540 51684 25596
rect 51684 25540 51740 25596
rect 51740 25540 51744 25596
rect 51680 25536 51744 25540
rect 51760 25596 51824 25600
rect 51760 25540 51764 25596
rect 51764 25540 51820 25596
rect 51820 25540 51824 25596
rect 51760 25536 51824 25540
rect 15400 25052 15464 25056
rect 15400 24996 15404 25052
rect 15404 24996 15460 25052
rect 15460 24996 15464 25052
rect 15400 24992 15464 24996
rect 15480 25052 15544 25056
rect 15480 24996 15484 25052
rect 15484 24996 15540 25052
rect 15540 24996 15544 25052
rect 15480 24992 15544 24996
rect 15560 25052 15624 25056
rect 15560 24996 15564 25052
rect 15564 24996 15620 25052
rect 15620 24996 15624 25052
rect 15560 24992 15624 24996
rect 15640 25052 15704 25056
rect 15640 24996 15644 25052
rect 15644 24996 15700 25052
rect 15700 24996 15704 25052
rect 15640 24992 15704 24996
rect 29848 25052 29912 25056
rect 29848 24996 29852 25052
rect 29852 24996 29908 25052
rect 29908 24996 29912 25052
rect 29848 24992 29912 24996
rect 29928 25052 29992 25056
rect 29928 24996 29932 25052
rect 29932 24996 29988 25052
rect 29988 24996 29992 25052
rect 29928 24992 29992 24996
rect 30008 25052 30072 25056
rect 30008 24996 30012 25052
rect 30012 24996 30068 25052
rect 30068 24996 30072 25052
rect 30008 24992 30072 24996
rect 30088 25052 30152 25056
rect 30088 24996 30092 25052
rect 30092 24996 30148 25052
rect 30148 24996 30152 25052
rect 30088 24992 30152 24996
rect 44296 25052 44360 25056
rect 44296 24996 44300 25052
rect 44300 24996 44356 25052
rect 44356 24996 44360 25052
rect 44296 24992 44360 24996
rect 44376 25052 44440 25056
rect 44376 24996 44380 25052
rect 44380 24996 44436 25052
rect 44436 24996 44440 25052
rect 44376 24992 44440 24996
rect 44456 25052 44520 25056
rect 44456 24996 44460 25052
rect 44460 24996 44516 25052
rect 44516 24996 44520 25052
rect 44456 24992 44520 24996
rect 44536 25052 44600 25056
rect 44536 24996 44540 25052
rect 44540 24996 44596 25052
rect 44596 24996 44600 25052
rect 44536 24992 44600 24996
rect 8176 24508 8240 24512
rect 8176 24452 8180 24508
rect 8180 24452 8236 24508
rect 8236 24452 8240 24508
rect 8176 24448 8240 24452
rect 8256 24508 8320 24512
rect 8256 24452 8260 24508
rect 8260 24452 8316 24508
rect 8316 24452 8320 24508
rect 8256 24448 8320 24452
rect 8336 24508 8400 24512
rect 8336 24452 8340 24508
rect 8340 24452 8396 24508
rect 8396 24452 8400 24508
rect 8336 24448 8400 24452
rect 8416 24508 8480 24512
rect 8416 24452 8420 24508
rect 8420 24452 8476 24508
rect 8476 24452 8480 24508
rect 8416 24448 8480 24452
rect 22624 24508 22688 24512
rect 22624 24452 22628 24508
rect 22628 24452 22684 24508
rect 22684 24452 22688 24508
rect 22624 24448 22688 24452
rect 22704 24508 22768 24512
rect 22704 24452 22708 24508
rect 22708 24452 22764 24508
rect 22764 24452 22768 24508
rect 22704 24448 22768 24452
rect 22784 24508 22848 24512
rect 22784 24452 22788 24508
rect 22788 24452 22844 24508
rect 22844 24452 22848 24508
rect 22784 24448 22848 24452
rect 22864 24508 22928 24512
rect 22864 24452 22868 24508
rect 22868 24452 22924 24508
rect 22924 24452 22928 24508
rect 22864 24448 22928 24452
rect 37072 24508 37136 24512
rect 37072 24452 37076 24508
rect 37076 24452 37132 24508
rect 37132 24452 37136 24508
rect 37072 24448 37136 24452
rect 37152 24508 37216 24512
rect 37152 24452 37156 24508
rect 37156 24452 37212 24508
rect 37212 24452 37216 24508
rect 37152 24448 37216 24452
rect 37232 24508 37296 24512
rect 37232 24452 37236 24508
rect 37236 24452 37292 24508
rect 37292 24452 37296 24508
rect 37232 24448 37296 24452
rect 37312 24508 37376 24512
rect 37312 24452 37316 24508
rect 37316 24452 37372 24508
rect 37372 24452 37376 24508
rect 37312 24448 37376 24452
rect 51520 24508 51584 24512
rect 51520 24452 51524 24508
rect 51524 24452 51580 24508
rect 51580 24452 51584 24508
rect 51520 24448 51584 24452
rect 51600 24508 51664 24512
rect 51600 24452 51604 24508
rect 51604 24452 51660 24508
rect 51660 24452 51664 24508
rect 51600 24448 51664 24452
rect 51680 24508 51744 24512
rect 51680 24452 51684 24508
rect 51684 24452 51740 24508
rect 51740 24452 51744 24508
rect 51680 24448 51744 24452
rect 51760 24508 51824 24512
rect 51760 24452 51764 24508
rect 51764 24452 51820 24508
rect 51820 24452 51824 24508
rect 51760 24448 51824 24452
rect 15400 23964 15464 23968
rect 15400 23908 15404 23964
rect 15404 23908 15460 23964
rect 15460 23908 15464 23964
rect 15400 23904 15464 23908
rect 15480 23964 15544 23968
rect 15480 23908 15484 23964
rect 15484 23908 15540 23964
rect 15540 23908 15544 23964
rect 15480 23904 15544 23908
rect 15560 23964 15624 23968
rect 15560 23908 15564 23964
rect 15564 23908 15620 23964
rect 15620 23908 15624 23964
rect 15560 23904 15624 23908
rect 15640 23964 15704 23968
rect 15640 23908 15644 23964
rect 15644 23908 15700 23964
rect 15700 23908 15704 23964
rect 15640 23904 15704 23908
rect 29848 23964 29912 23968
rect 29848 23908 29852 23964
rect 29852 23908 29908 23964
rect 29908 23908 29912 23964
rect 29848 23904 29912 23908
rect 29928 23964 29992 23968
rect 29928 23908 29932 23964
rect 29932 23908 29988 23964
rect 29988 23908 29992 23964
rect 29928 23904 29992 23908
rect 30008 23964 30072 23968
rect 30008 23908 30012 23964
rect 30012 23908 30068 23964
rect 30068 23908 30072 23964
rect 30008 23904 30072 23908
rect 30088 23964 30152 23968
rect 30088 23908 30092 23964
rect 30092 23908 30148 23964
rect 30148 23908 30152 23964
rect 30088 23904 30152 23908
rect 44296 23964 44360 23968
rect 44296 23908 44300 23964
rect 44300 23908 44356 23964
rect 44356 23908 44360 23964
rect 44296 23904 44360 23908
rect 44376 23964 44440 23968
rect 44376 23908 44380 23964
rect 44380 23908 44436 23964
rect 44436 23908 44440 23964
rect 44376 23904 44440 23908
rect 44456 23964 44520 23968
rect 44456 23908 44460 23964
rect 44460 23908 44516 23964
rect 44516 23908 44520 23964
rect 44456 23904 44520 23908
rect 44536 23964 44600 23968
rect 44536 23908 44540 23964
rect 44540 23908 44596 23964
rect 44596 23908 44600 23964
rect 44536 23904 44600 23908
rect 8176 23420 8240 23424
rect 8176 23364 8180 23420
rect 8180 23364 8236 23420
rect 8236 23364 8240 23420
rect 8176 23360 8240 23364
rect 8256 23420 8320 23424
rect 8256 23364 8260 23420
rect 8260 23364 8316 23420
rect 8316 23364 8320 23420
rect 8256 23360 8320 23364
rect 8336 23420 8400 23424
rect 8336 23364 8340 23420
rect 8340 23364 8396 23420
rect 8396 23364 8400 23420
rect 8336 23360 8400 23364
rect 8416 23420 8480 23424
rect 8416 23364 8420 23420
rect 8420 23364 8476 23420
rect 8476 23364 8480 23420
rect 8416 23360 8480 23364
rect 22624 23420 22688 23424
rect 22624 23364 22628 23420
rect 22628 23364 22684 23420
rect 22684 23364 22688 23420
rect 22624 23360 22688 23364
rect 22704 23420 22768 23424
rect 22704 23364 22708 23420
rect 22708 23364 22764 23420
rect 22764 23364 22768 23420
rect 22704 23360 22768 23364
rect 22784 23420 22848 23424
rect 22784 23364 22788 23420
rect 22788 23364 22844 23420
rect 22844 23364 22848 23420
rect 22784 23360 22848 23364
rect 22864 23420 22928 23424
rect 22864 23364 22868 23420
rect 22868 23364 22924 23420
rect 22924 23364 22928 23420
rect 22864 23360 22928 23364
rect 37072 23420 37136 23424
rect 37072 23364 37076 23420
rect 37076 23364 37132 23420
rect 37132 23364 37136 23420
rect 37072 23360 37136 23364
rect 37152 23420 37216 23424
rect 37152 23364 37156 23420
rect 37156 23364 37212 23420
rect 37212 23364 37216 23420
rect 37152 23360 37216 23364
rect 37232 23420 37296 23424
rect 37232 23364 37236 23420
rect 37236 23364 37292 23420
rect 37292 23364 37296 23420
rect 37232 23360 37296 23364
rect 37312 23420 37376 23424
rect 37312 23364 37316 23420
rect 37316 23364 37372 23420
rect 37372 23364 37376 23420
rect 37312 23360 37376 23364
rect 51520 23420 51584 23424
rect 51520 23364 51524 23420
rect 51524 23364 51580 23420
rect 51580 23364 51584 23420
rect 51520 23360 51584 23364
rect 51600 23420 51664 23424
rect 51600 23364 51604 23420
rect 51604 23364 51660 23420
rect 51660 23364 51664 23420
rect 51600 23360 51664 23364
rect 51680 23420 51744 23424
rect 51680 23364 51684 23420
rect 51684 23364 51740 23420
rect 51740 23364 51744 23420
rect 51680 23360 51744 23364
rect 51760 23420 51824 23424
rect 51760 23364 51764 23420
rect 51764 23364 51820 23420
rect 51820 23364 51824 23420
rect 51760 23360 51824 23364
rect 15400 22876 15464 22880
rect 15400 22820 15404 22876
rect 15404 22820 15460 22876
rect 15460 22820 15464 22876
rect 15400 22816 15464 22820
rect 15480 22876 15544 22880
rect 15480 22820 15484 22876
rect 15484 22820 15540 22876
rect 15540 22820 15544 22876
rect 15480 22816 15544 22820
rect 15560 22876 15624 22880
rect 15560 22820 15564 22876
rect 15564 22820 15620 22876
rect 15620 22820 15624 22876
rect 15560 22816 15624 22820
rect 15640 22876 15704 22880
rect 15640 22820 15644 22876
rect 15644 22820 15700 22876
rect 15700 22820 15704 22876
rect 15640 22816 15704 22820
rect 29848 22876 29912 22880
rect 29848 22820 29852 22876
rect 29852 22820 29908 22876
rect 29908 22820 29912 22876
rect 29848 22816 29912 22820
rect 29928 22876 29992 22880
rect 29928 22820 29932 22876
rect 29932 22820 29988 22876
rect 29988 22820 29992 22876
rect 29928 22816 29992 22820
rect 30008 22876 30072 22880
rect 30008 22820 30012 22876
rect 30012 22820 30068 22876
rect 30068 22820 30072 22876
rect 30008 22816 30072 22820
rect 30088 22876 30152 22880
rect 30088 22820 30092 22876
rect 30092 22820 30148 22876
rect 30148 22820 30152 22876
rect 30088 22816 30152 22820
rect 44296 22876 44360 22880
rect 44296 22820 44300 22876
rect 44300 22820 44356 22876
rect 44356 22820 44360 22876
rect 44296 22816 44360 22820
rect 44376 22876 44440 22880
rect 44376 22820 44380 22876
rect 44380 22820 44436 22876
rect 44436 22820 44440 22876
rect 44376 22816 44440 22820
rect 44456 22876 44520 22880
rect 44456 22820 44460 22876
rect 44460 22820 44516 22876
rect 44516 22820 44520 22876
rect 44456 22816 44520 22820
rect 44536 22876 44600 22880
rect 44536 22820 44540 22876
rect 44540 22820 44596 22876
rect 44596 22820 44600 22876
rect 44536 22816 44600 22820
rect 8176 22332 8240 22336
rect 8176 22276 8180 22332
rect 8180 22276 8236 22332
rect 8236 22276 8240 22332
rect 8176 22272 8240 22276
rect 8256 22332 8320 22336
rect 8256 22276 8260 22332
rect 8260 22276 8316 22332
rect 8316 22276 8320 22332
rect 8256 22272 8320 22276
rect 8336 22332 8400 22336
rect 8336 22276 8340 22332
rect 8340 22276 8396 22332
rect 8396 22276 8400 22332
rect 8336 22272 8400 22276
rect 8416 22332 8480 22336
rect 8416 22276 8420 22332
rect 8420 22276 8476 22332
rect 8476 22276 8480 22332
rect 8416 22272 8480 22276
rect 22624 22332 22688 22336
rect 22624 22276 22628 22332
rect 22628 22276 22684 22332
rect 22684 22276 22688 22332
rect 22624 22272 22688 22276
rect 22704 22332 22768 22336
rect 22704 22276 22708 22332
rect 22708 22276 22764 22332
rect 22764 22276 22768 22332
rect 22704 22272 22768 22276
rect 22784 22332 22848 22336
rect 22784 22276 22788 22332
rect 22788 22276 22844 22332
rect 22844 22276 22848 22332
rect 22784 22272 22848 22276
rect 22864 22332 22928 22336
rect 22864 22276 22868 22332
rect 22868 22276 22924 22332
rect 22924 22276 22928 22332
rect 22864 22272 22928 22276
rect 37072 22332 37136 22336
rect 37072 22276 37076 22332
rect 37076 22276 37132 22332
rect 37132 22276 37136 22332
rect 37072 22272 37136 22276
rect 37152 22332 37216 22336
rect 37152 22276 37156 22332
rect 37156 22276 37212 22332
rect 37212 22276 37216 22332
rect 37152 22272 37216 22276
rect 37232 22332 37296 22336
rect 37232 22276 37236 22332
rect 37236 22276 37292 22332
rect 37292 22276 37296 22332
rect 37232 22272 37296 22276
rect 37312 22332 37376 22336
rect 37312 22276 37316 22332
rect 37316 22276 37372 22332
rect 37372 22276 37376 22332
rect 37312 22272 37376 22276
rect 51520 22332 51584 22336
rect 51520 22276 51524 22332
rect 51524 22276 51580 22332
rect 51580 22276 51584 22332
rect 51520 22272 51584 22276
rect 51600 22332 51664 22336
rect 51600 22276 51604 22332
rect 51604 22276 51660 22332
rect 51660 22276 51664 22332
rect 51600 22272 51664 22276
rect 51680 22332 51744 22336
rect 51680 22276 51684 22332
rect 51684 22276 51740 22332
rect 51740 22276 51744 22332
rect 51680 22272 51744 22276
rect 51760 22332 51824 22336
rect 51760 22276 51764 22332
rect 51764 22276 51820 22332
rect 51820 22276 51824 22332
rect 51760 22272 51824 22276
rect 15400 21788 15464 21792
rect 15400 21732 15404 21788
rect 15404 21732 15460 21788
rect 15460 21732 15464 21788
rect 15400 21728 15464 21732
rect 15480 21788 15544 21792
rect 15480 21732 15484 21788
rect 15484 21732 15540 21788
rect 15540 21732 15544 21788
rect 15480 21728 15544 21732
rect 15560 21788 15624 21792
rect 15560 21732 15564 21788
rect 15564 21732 15620 21788
rect 15620 21732 15624 21788
rect 15560 21728 15624 21732
rect 15640 21788 15704 21792
rect 15640 21732 15644 21788
rect 15644 21732 15700 21788
rect 15700 21732 15704 21788
rect 15640 21728 15704 21732
rect 29848 21788 29912 21792
rect 29848 21732 29852 21788
rect 29852 21732 29908 21788
rect 29908 21732 29912 21788
rect 29848 21728 29912 21732
rect 29928 21788 29992 21792
rect 29928 21732 29932 21788
rect 29932 21732 29988 21788
rect 29988 21732 29992 21788
rect 29928 21728 29992 21732
rect 30008 21788 30072 21792
rect 30008 21732 30012 21788
rect 30012 21732 30068 21788
rect 30068 21732 30072 21788
rect 30008 21728 30072 21732
rect 30088 21788 30152 21792
rect 30088 21732 30092 21788
rect 30092 21732 30148 21788
rect 30148 21732 30152 21788
rect 30088 21728 30152 21732
rect 44296 21788 44360 21792
rect 44296 21732 44300 21788
rect 44300 21732 44356 21788
rect 44356 21732 44360 21788
rect 44296 21728 44360 21732
rect 44376 21788 44440 21792
rect 44376 21732 44380 21788
rect 44380 21732 44436 21788
rect 44436 21732 44440 21788
rect 44376 21728 44440 21732
rect 44456 21788 44520 21792
rect 44456 21732 44460 21788
rect 44460 21732 44516 21788
rect 44516 21732 44520 21788
rect 44456 21728 44520 21732
rect 44536 21788 44600 21792
rect 44536 21732 44540 21788
rect 44540 21732 44596 21788
rect 44596 21732 44600 21788
rect 44536 21728 44600 21732
rect 8176 21244 8240 21248
rect 8176 21188 8180 21244
rect 8180 21188 8236 21244
rect 8236 21188 8240 21244
rect 8176 21184 8240 21188
rect 8256 21244 8320 21248
rect 8256 21188 8260 21244
rect 8260 21188 8316 21244
rect 8316 21188 8320 21244
rect 8256 21184 8320 21188
rect 8336 21244 8400 21248
rect 8336 21188 8340 21244
rect 8340 21188 8396 21244
rect 8396 21188 8400 21244
rect 8336 21184 8400 21188
rect 8416 21244 8480 21248
rect 8416 21188 8420 21244
rect 8420 21188 8476 21244
rect 8476 21188 8480 21244
rect 8416 21184 8480 21188
rect 22624 21244 22688 21248
rect 22624 21188 22628 21244
rect 22628 21188 22684 21244
rect 22684 21188 22688 21244
rect 22624 21184 22688 21188
rect 22704 21244 22768 21248
rect 22704 21188 22708 21244
rect 22708 21188 22764 21244
rect 22764 21188 22768 21244
rect 22704 21184 22768 21188
rect 22784 21244 22848 21248
rect 22784 21188 22788 21244
rect 22788 21188 22844 21244
rect 22844 21188 22848 21244
rect 22784 21184 22848 21188
rect 22864 21244 22928 21248
rect 22864 21188 22868 21244
rect 22868 21188 22924 21244
rect 22924 21188 22928 21244
rect 22864 21184 22928 21188
rect 37072 21244 37136 21248
rect 37072 21188 37076 21244
rect 37076 21188 37132 21244
rect 37132 21188 37136 21244
rect 37072 21184 37136 21188
rect 37152 21244 37216 21248
rect 37152 21188 37156 21244
rect 37156 21188 37212 21244
rect 37212 21188 37216 21244
rect 37152 21184 37216 21188
rect 37232 21244 37296 21248
rect 37232 21188 37236 21244
rect 37236 21188 37292 21244
rect 37292 21188 37296 21244
rect 37232 21184 37296 21188
rect 37312 21244 37376 21248
rect 37312 21188 37316 21244
rect 37316 21188 37372 21244
rect 37372 21188 37376 21244
rect 37312 21184 37376 21188
rect 51520 21244 51584 21248
rect 51520 21188 51524 21244
rect 51524 21188 51580 21244
rect 51580 21188 51584 21244
rect 51520 21184 51584 21188
rect 51600 21244 51664 21248
rect 51600 21188 51604 21244
rect 51604 21188 51660 21244
rect 51660 21188 51664 21244
rect 51600 21184 51664 21188
rect 51680 21244 51744 21248
rect 51680 21188 51684 21244
rect 51684 21188 51740 21244
rect 51740 21188 51744 21244
rect 51680 21184 51744 21188
rect 51760 21244 51824 21248
rect 51760 21188 51764 21244
rect 51764 21188 51820 21244
rect 51820 21188 51824 21244
rect 51760 21184 51824 21188
rect 15400 20700 15464 20704
rect 15400 20644 15404 20700
rect 15404 20644 15460 20700
rect 15460 20644 15464 20700
rect 15400 20640 15464 20644
rect 15480 20700 15544 20704
rect 15480 20644 15484 20700
rect 15484 20644 15540 20700
rect 15540 20644 15544 20700
rect 15480 20640 15544 20644
rect 15560 20700 15624 20704
rect 15560 20644 15564 20700
rect 15564 20644 15620 20700
rect 15620 20644 15624 20700
rect 15560 20640 15624 20644
rect 15640 20700 15704 20704
rect 15640 20644 15644 20700
rect 15644 20644 15700 20700
rect 15700 20644 15704 20700
rect 15640 20640 15704 20644
rect 29848 20700 29912 20704
rect 29848 20644 29852 20700
rect 29852 20644 29908 20700
rect 29908 20644 29912 20700
rect 29848 20640 29912 20644
rect 29928 20700 29992 20704
rect 29928 20644 29932 20700
rect 29932 20644 29988 20700
rect 29988 20644 29992 20700
rect 29928 20640 29992 20644
rect 30008 20700 30072 20704
rect 30008 20644 30012 20700
rect 30012 20644 30068 20700
rect 30068 20644 30072 20700
rect 30008 20640 30072 20644
rect 30088 20700 30152 20704
rect 30088 20644 30092 20700
rect 30092 20644 30148 20700
rect 30148 20644 30152 20700
rect 30088 20640 30152 20644
rect 44296 20700 44360 20704
rect 44296 20644 44300 20700
rect 44300 20644 44356 20700
rect 44356 20644 44360 20700
rect 44296 20640 44360 20644
rect 44376 20700 44440 20704
rect 44376 20644 44380 20700
rect 44380 20644 44436 20700
rect 44436 20644 44440 20700
rect 44376 20640 44440 20644
rect 44456 20700 44520 20704
rect 44456 20644 44460 20700
rect 44460 20644 44516 20700
rect 44516 20644 44520 20700
rect 44456 20640 44520 20644
rect 44536 20700 44600 20704
rect 44536 20644 44540 20700
rect 44540 20644 44596 20700
rect 44596 20644 44600 20700
rect 44536 20640 44600 20644
rect 8176 20156 8240 20160
rect 8176 20100 8180 20156
rect 8180 20100 8236 20156
rect 8236 20100 8240 20156
rect 8176 20096 8240 20100
rect 8256 20156 8320 20160
rect 8256 20100 8260 20156
rect 8260 20100 8316 20156
rect 8316 20100 8320 20156
rect 8256 20096 8320 20100
rect 8336 20156 8400 20160
rect 8336 20100 8340 20156
rect 8340 20100 8396 20156
rect 8396 20100 8400 20156
rect 8336 20096 8400 20100
rect 8416 20156 8480 20160
rect 8416 20100 8420 20156
rect 8420 20100 8476 20156
rect 8476 20100 8480 20156
rect 8416 20096 8480 20100
rect 22624 20156 22688 20160
rect 22624 20100 22628 20156
rect 22628 20100 22684 20156
rect 22684 20100 22688 20156
rect 22624 20096 22688 20100
rect 22704 20156 22768 20160
rect 22704 20100 22708 20156
rect 22708 20100 22764 20156
rect 22764 20100 22768 20156
rect 22704 20096 22768 20100
rect 22784 20156 22848 20160
rect 22784 20100 22788 20156
rect 22788 20100 22844 20156
rect 22844 20100 22848 20156
rect 22784 20096 22848 20100
rect 22864 20156 22928 20160
rect 22864 20100 22868 20156
rect 22868 20100 22924 20156
rect 22924 20100 22928 20156
rect 22864 20096 22928 20100
rect 37072 20156 37136 20160
rect 37072 20100 37076 20156
rect 37076 20100 37132 20156
rect 37132 20100 37136 20156
rect 37072 20096 37136 20100
rect 37152 20156 37216 20160
rect 37152 20100 37156 20156
rect 37156 20100 37212 20156
rect 37212 20100 37216 20156
rect 37152 20096 37216 20100
rect 37232 20156 37296 20160
rect 37232 20100 37236 20156
rect 37236 20100 37292 20156
rect 37292 20100 37296 20156
rect 37232 20096 37296 20100
rect 37312 20156 37376 20160
rect 37312 20100 37316 20156
rect 37316 20100 37372 20156
rect 37372 20100 37376 20156
rect 37312 20096 37376 20100
rect 51520 20156 51584 20160
rect 51520 20100 51524 20156
rect 51524 20100 51580 20156
rect 51580 20100 51584 20156
rect 51520 20096 51584 20100
rect 51600 20156 51664 20160
rect 51600 20100 51604 20156
rect 51604 20100 51660 20156
rect 51660 20100 51664 20156
rect 51600 20096 51664 20100
rect 51680 20156 51744 20160
rect 51680 20100 51684 20156
rect 51684 20100 51740 20156
rect 51740 20100 51744 20156
rect 51680 20096 51744 20100
rect 51760 20156 51824 20160
rect 51760 20100 51764 20156
rect 51764 20100 51820 20156
rect 51820 20100 51824 20156
rect 51760 20096 51824 20100
rect 15400 19612 15464 19616
rect 15400 19556 15404 19612
rect 15404 19556 15460 19612
rect 15460 19556 15464 19612
rect 15400 19552 15464 19556
rect 15480 19612 15544 19616
rect 15480 19556 15484 19612
rect 15484 19556 15540 19612
rect 15540 19556 15544 19612
rect 15480 19552 15544 19556
rect 15560 19612 15624 19616
rect 15560 19556 15564 19612
rect 15564 19556 15620 19612
rect 15620 19556 15624 19612
rect 15560 19552 15624 19556
rect 15640 19612 15704 19616
rect 15640 19556 15644 19612
rect 15644 19556 15700 19612
rect 15700 19556 15704 19612
rect 15640 19552 15704 19556
rect 29848 19612 29912 19616
rect 29848 19556 29852 19612
rect 29852 19556 29908 19612
rect 29908 19556 29912 19612
rect 29848 19552 29912 19556
rect 29928 19612 29992 19616
rect 29928 19556 29932 19612
rect 29932 19556 29988 19612
rect 29988 19556 29992 19612
rect 29928 19552 29992 19556
rect 30008 19612 30072 19616
rect 30008 19556 30012 19612
rect 30012 19556 30068 19612
rect 30068 19556 30072 19612
rect 30008 19552 30072 19556
rect 30088 19612 30152 19616
rect 30088 19556 30092 19612
rect 30092 19556 30148 19612
rect 30148 19556 30152 19612
rect 30088 19552 30152 19556
rect 44296 19612 44360 19616
rect 44296 19556 44300 19612
rect 44300 19556 44356 19612
rect 44356 19556 44360 19612
rect 44296 19552 44360 19556
rect 44376 19612 44440 19616
rect 44376 19556 44380 19612
rect 44380 19556 44436 19612
rect 44436 19556 44440 19612
rect 44376 19552 44440 19556
rect 44456 19612 44520 19616
rect 44456 19556 44460 19612
rect 44460 19556 44516 19612
rect 44516 19556 44520 19612
rect 44456 19552 44520 19556
rect 44536 19612 44600 19616
rect 44536 19556 44540 19612
rect 44540 19556 44596 19612
rect 44596 19556 44600 19612
rect 44536 19552 44600 19556
rect 8176 19068 8240 19072
rect 8176 19012 8180 19068
rect 8180 19012 8236 19068
rect 8236 19012 8240 19068
rect 8176 19008 8240 19012
rect 8256 19068 8320 19072
rect 8256 19012 8260 19068
rect 8260 19012 8316 19068
rect 8316 19012 8320 19068
rect 8256 19008 8320 19012
rect 8336 19068 8400 19072
rect 8336 19012 8340 19068
rect 8340 19012 8396 19068
rect 8396 19012 8400 19068
rect 8336 19008 8400 19012
rect 8416 19068 8480 19072
rect 8416 19012 8420 19068
rect 8420 19012 8476 19068
rect 8476 19012 8480 19068
rect 8416 19008 8480 19012
rect 22624 19068 22688 19072
rect 22624 19012 22628 19068
rect 22628 19012 22684 19068
rect 22684 19012 22688 19068
rect 22624 19008 22688 19012
rect 22704 19068 22768 19072
rect 22704 19012 22708 19068
rect 22708 19012 22764 19068
rect 22764 19012 22768 19068
rect 22704 19008 22768 19012
rect 22784 19068 22848 19072
rect 22784 19012 22788 19068
rect 22788 19012 22844 19068
rect 22844 19012 22848 19068
rect 22784 19008 22848 19012
rect 22864 19068 22928 19072
rect 22864 19012 22868 19068
rect 22868 19012 22924 19068
rect 22924 19012 22928 19068
rect 22864 19008 22928 19012
rect 37072 19068 37136 19072
rect 37072 19012 37076 19068
rect 37076 19012 37132 19068
rect 37132 19012 37136 19068
rect 37072 19008 37136 19012
rect 37152 19068 37216 19072
rect 37152 19012 37156 19068
rect 37156 19012 37212 19068
rect 37212 19012 37216 19068
rect 37152 19008 37216 19012
rect 37232 19068 37296 19072
rect 37232 19012 37236 19068
rect 37236 19012 37292 19068
rect 37292 19012 37296 19068
rect 37232 19008 37296 19012
rect 37312 19068 37376 19072
rect 37312 19012 37316 19068
rect 37316 19012 37372 19068
rect 37372 19012 37376 19068
rect 37312 19008 37376 19012
rect 51520 19068 51584 19072
rect 51520 19012 51524 19068
rect 51524 19012 51580 19068
rect 51580 19012 51584 19068
rect 51520 19008 51584 19012
rect 51600 19068 51664 19072
rect 51600 19012 51604 19068
rect 51604 19012 51660 19068
rect 51660 19012 51664 19068
rect 51600 19008 51664 19012
rect 51680 19068 51744 19072
rect 51680 19012 51684 19068
rect 51684 19012 51740 19068
rect 51740 19012 51744 19068
rect 51680 19008 51744 19012
rect 51760 19068 51824 19072
rect 51760 19012 51764 19068
rect 51764 19012 51820 19068
rect 51820 19012 51824 19068
rect 51760 19008 51824 19012
rect 15400 18524 15464 18528
rect 15400 18468 15404 18524
rect 15404 18468 15460 18524
rect 15460 18468 15464 18524
rect 15400 18464 15464 18468
rect 15480 18524 15544 18528
rect 15480 18468 15484 18524
rect 15484 18468 15540 18524
rect 15540 18468 15544 18524
rect 15480 18464 15544 18468
rect 15560 18524 15624 18528
rect 15560 18468 15564 18524
rect 15564 18468 15620 18524
rect 15620 18468 15624 18524
rect 15560 18464 15624 18468
rect 15640 18524 15704 18528
rect 15640 18468 15644 18524
rect 15644 18468 15700 18524
rect 15700 18468 15704 18524
rect 15640 18464 15704 18468
rect 29848 18524 29912 18528
rect 29848 18468 29852 18524
rect 29852 18468 29908 18524
rect 29908 18468 29912 18524
rect 29848 18464 29912 18468
rect 29928 18524 29992 18528
rect 29928 18468 29932 18524
rect 29932 18468 29988 18524
rect 29988 18468 29992 18524
rect 29928 18464 29992 18468
rect 30008 18524 30072 18528
rect 30008 18468 30012 18524
rect 30012 18468 30068 18524
rect 30068 18468 30072 18524
rect 30008 18464 30072 18468
rect 30088 18524 30152 18528
rect 30088 18468 30092 18524
rect 30092 18468 30148 18524
rect 30148 18468 30152 18524
rect 30088 18464 30152 18468
rect 44296 18524 44360 18528
rect 44296 18468 44300 18524
rect 44300 18468 44356 18524
rect 44356 18468 44360 18524
rect 44296 18464 44360 18468
rect 44376 18524 44440 18528
rect 44376 18468 44380 18524
rect 44380 18468 44436 18524
rect 44436 18468 44440 18524
rect 44376 18464 44440 18468
rect 44456 18524 44520 18528
rect 44456 18468 44460 18524
rect 44460 18468 44516 18524
rect 44516 18468 44520 18524
rect 44456 18464 44520 18468
rect 44536 18524 44600 18528
rect 44536 18468 44540 18524
rect 44540 18468 44596 18524
rect 44596 18468 44600 18524
rect 44536 18464 44600 18468
rect 8176 17980 8240 17984
rect 8176 17924 8180 17980
rect 8180 17924 8236 17980
rect 8236 17924 8240 17980
rect 8176 17920 8240 17924
rect 8256 17980 8320 17984
rect 8256 17924 8260 17980
rect 8260 17924 8316 17980
rect 8316 17924 8320 17980
rect 8256 17920 8320 17924
rect 8336 17980 8400 17984
rect 8336 17924 8340 17980
rect 8340 17924 8396 17980
rect 8396 17924 8400 17980
rect 8336 17920 8400 17924
rect 8416 17980 8480 17984
rect 8416 17924 8420 17980
rect 8420 17924 8476 17980
rect 8476 17924 8480 17980
rect 8416 17920 8480 17924
rect 22624 17980 22688 17984
rect 22624 17924 22628 17980
rect 22628 17924 22684 17980
rect 22684 17924 22688 17980
rect 22624 17920 22688 17924
rect 22704 17980 22768 17984
rect 22704 17924 22708 17980
rect 22708 17924 22764 17980
rect 22764 17924 22768 17980
rect 22704 17920 22768 17924
rect 22784 17980 22848 17984
rect 22784 17924 22788 17980
rect 22788 17924 22844 17980
rect 22844 17924 22848 17980
rect 22784 17920 22848 17924
rect 22864 17980 22928 17984
rect 22864 17924 22868 17980
rect 22868 17924 22924 17980
rect 22924 17924 22928 17980
rect 22864 17920 22928 17924
rect 37072 17980 37136 17984
rect 37072 17924 37076 17980
rect 37076 17924 37132 17980
rect 37132 17924 37136 17980
rect 37072 17920 37136 17924
rect 37152 17980 37216 17984
rect 37152 17924 37156 17980
rect 37156 17924 37212 17980
rect 37212 17924 37216 17980
rect 37152 17920 37216 17924
rect 37232 17980 37296 17984
rect 37232 17924 37236 17980
rect 37236 17924 37292 17980
rect 37292 17924 37296 17980
rect 37232 17920 37296 17924
rect 37312 17980 37376 17984
rect 37312 17924 37316 17980
rect 37316 17924 37372 17980
rect 37372 17924 37376 17980
rect 37312 17920 37376 17924
rect 51520 17980 51584 17984
rect 51520 17924 51524 17980
rect 51524 17924 51580 17980
rect 51580 17924 51584 17980
rect 51520 17920 51584 17924
rect 51600 17980 51664 17984
rect 51600 17924 51604 17980
rect 51604 17924 51660 17980
rect 51660 17924 51664 17980
rect 51600 17920 51664 17924
rect 51680 17980 51744 17984
rect 51680 17924 51684 17980
rect 51684 17924 51740 17980
rect 51740 17924 51744 17980
rect 51680 17920 51744 17924
rect 51760 17980 51824 17984
rect 51760 17924 51764 17980
rect 51764 17924 51820 17980
rect 51820 17924 51824 17980
rect 51760 17920 51824 17924
rect 15400 17436 15464 17440
rect 15400 17380 15404 17436
rect 15404 17380 15460 17436
rect 15460 17380 15464 17436
rect 15400 17376 15464 17380
rect 15480 17436 15544 17440
rect 15480 17380 15484 17436
rect 15484 17380 15540 17436
rect 15540 17380 15544 17436
rect 15480 17376 15544 17380
rect 15560 17436 15624 17440
rect 15560 17380 15564 17436
rect 15564 17380 15620 17436
rect 15620 17380 15624 17436
rect 15560 17376 15624 17380
rect 15640 17436 15704 17440
rect 15640 17380 15644 17436
rect 15644 17380 15700 17436
rect 15700 17380 15704 17436
rect 15640 17376 15704 17380
rect 29848 17436 29912 17440
rect 29848 17380 29852 17436
rect 29852 17380 29908 17436
rect 29908 17380 29912 17436
rect 29848 17376 29912 17380
rect 29928 17436 29992 17440
rect 29928 17380 29932 17436
rect 29932 17380 29988 17436
rect 29988 17380 29992 17436
rect 29928 17376 29992 17380
rect 30008 17436 30072 17440
rect 30008 17380 30012 17436
rect 30012 17380 30068 17436
rect 30068 17380 30072 17436
rect 30008 17376 30072 17380
rect 30088 17436 30152 17440
rect 30088 17380 30092 17436
rect 30092 17380 30148 17436
rect 30148 17380 30152 17436
rect 30088 17376 30152 17380
rect 44296 17436 44360 17440
rect 44296 17380 44300 17436
rect 44300 17380 44356 17436
rect 44356 17380 44360 17436
rect 44296 17376 44360 17380
rect 44376 17436 44440 17440
rect 44376 17380 44380 17436
rect 44380 17380 44436 17436
rect 44436 17380 44440 17436
rect 44376 17376 44440 17380
rect 44456 17436 44520 17440
rect 44456 17380 44460 17436
rect 44460 17380 44516 17436
rect 44516 17380 44520 17436
rect 44456 17376 44520 17380
rect 44536 17436 44600 17440
rect 44536 17380 44540 17436
rect 44540 17380 44596 17436
rect 44596 17380 44600 17436
rect 44536 17376 44600 17380
rect 8176 16892 8240 16896
rect 8176 16836 8180 16892
rect 8180 16836 8236 16892
rect 8236 16836 8240 16892
rect 8176 16832 8240 16836
rect 8256 16892 8320 16896
rect 8256 16836 8260 16892
rect 8260 16836 8316 16892
rect 8316 16836 8320 16892
rect 8256 16832 8320 16836
rect 8336 16892 8400 16896
rect 8336 16836 8340 16892
rect 8340 16836 8396 16892
rect 8396 16836 8400 16892
rect 8336 16832 8400 16836
rect 8416 16892 8480 16896
rect 8416 16836 8420 16892
rect 8420 16836 8476 16892
rect 8476 16836 8480 16892
rect 8416 16832 8480 16836
rect 22624 16892 22688 16896
rect 22624 16836 22628 16892
rect 22628 16836 22684 16892
rect 22684 16836 22688 16892
rect 22624 16832 22688 16836
rect 22704 16892 22768 16896
rect 22704 16836 22708 16892
rect 22708 16836 22764 16892
rect 22764 16836 22768 16892
rect 22704 16832 22768 16836
rect 22784 16892 22848 16896
rect 22784 16836 22788 16892
rect 22788 16836 22844 16892
rect 22844 16836 22848 16892
rect 22784 16832 22848 16836
rect 22864 16892 22928 16896
rect 22864 16836 22868 16892
rect 22868 16836 22924 16892
rect 22924 16836 22928 16892
rect 22864 16832 22928 16836
rect 37072 16892 37136 16896
rect 37072 16836 37076 16892
rect 37076 16836 37132 16892
rect 37132 16836 37136 16892
rect 37072 16832 37136 16836
rect 37152 16892 37216 16896
rect 37152 16836 37156 16892
rect 37156 16836 37212 16892
rect 37212 16836 37216 16892
rect 37152 16832 37216 16836
rect 37232 16892 37296 16896
rect 37232 16836 37236 16892
rect 37236 16836 37292 16892
rect 37292 16836 37296 16892
rect 37232 16832 37296 16836
rect 37312 16892 37376 16896
rect 37312 16836 37316 16892
rect 37316 16836 37372 16892
rect 37372 16836 37376 16892
rect 37312 16832 37376 16836
rect 51520 16892 51584 16896
rect 51520 16836 51524 16892
rect 51524 16836 51580 16892
rect 51580 16836 51584 16892
rect 51520 16832 51584 16836
rect 51600 16892 51664 16896
rect 51600 16836 51604 16892
rect 51604 16836 51660 16892
rect 51660 16836 51664 16892
rect 51600 16832 51664 16836
rect 51680 16892 51744 16896
rect 51680 16836 51684 16892
rect 51684 16836 51740 16892
rect 51740 16836 51744 16892
rect 51680 16832 51744 16836
rect 51760 16892 51824 16896
rect 51760 16836 51764 16892
rect 51764 16836 51820 16892
rect 51820 16836 51824 16892
rect 51760 16832 51824 16836
rect 15400 16348 15464 16352
rect 15400 16292 15404 16348
rect 15404 16292 15460 16348
rect 15460 16292 15464 16348
rect 15400 16288 15464 16292
rect 15480 16348 15544 16352
rect 15480 16292 15484 16348
rect 15484 16292 15540 16348
rect 15540 16292 15544 16348
rect 15480 16288 15544 16292
rect 15560 16348 15624 16352
rect 15560 16292 15564 16348
rect 15564 16292 15620 16348
rect 15620 16292 15624 16348
rect 15560 16288 15624 16292
rect 15640 16348 15704 16352
rect 15640 16292 15644 16348
rect 15644 16292 15700 16348
rect 15700 16292 15704 16348
rect 15640 16288 15704 16292
rect 29848 16348 29912 16352
rect 29848 16292 29852 16348
rect 29852 16292 29908 16348
rect 29908 16292 29912 16348
rect 29848 16288 29912 16292
rect 29928 16348 29992 16352
rect 29928 16292 29932 16348
rect 29932 16292 29988 16348
rect 29988 16292 29992 16348
rect 29928 16288 29992 16292
rect 30008 16348 30072 16352
rect 30008 16292 30012 16348
rect 30012 16292 30068 16348
rect 30068 16292 30072 16348
rect 30008 16288 30072 16292
rect 30088 16348 30152 16352
rect 30088 16292 30092 16348
rect 30092 16292 30148 16348
rect 30148 16292 30152 16348
rect 30088 16288 30152 16292
rect 44296 16348 44360 16352
rect 44296 16292 44300 16348
rect 44300 16292 44356 16348
rect 44356 16292 44360 16348
rect 44296 16288 44360 16292
rect 44376 16348 44440 16352
rect 44376 16292 44380 16348
rect 44380 16292 44436 16348
rect 44436 16292 44440 16348
rect 44376 16288 44440 16292
rect 44456 16348 44520 16352
rect 44456 16292 44460 16348
rect 44460 16292 44516 16348
rect 44516 16292 44520 16348
rect 44456 16288 44520 16292
rect 44536 16348 44600 16352
rect 44536 16292 44540 16348
rect 44540 16292 44596 16348
rect 44596 16292 44600 16348
rect 44536 16288 44600 16292
rect 8176 15804 8240 15808
rect 8176 15748 8180 15804
rect 8180 15748 8236 15804
rect 8236 15748 8240 15804
rect 8176 15744 8240 15748
rect 8256 15804 8320 15808
rect 8256 15748 8260 15804
rect 8260 15748 8316 15804
rect 8316 15748 8320 15804
rect 8256 15744 8320 15748
rect 8336 15804 8400 15808
rect 8336 15748 8340 15804
rect 8340 15748 8396 15804
rect 8396 15748 8400 15804
rect 8336 15744 8400 15748
rect 8416 15804 8480 15808
rect 8416 15748 8420 15804
rect 8420 15748 8476 15804
rect 8476 15748 8480 15804
rect 8416 15744 8480 15748
rect 22624 15804 22688 15808
rect 22624 15748 22628 15804
rect 22628 15748 22684 15804
rect 22684 15748 22688 15804
rect 22624 15744 22688 15748
rect 22704 15804 22768 15808
rect 22704 15748 22708 15804
rect 22708 15748 22764 15804
rect 22764 15748 22768 15804
rect 22704 15744 22768 15748
rect 22784 15804 22848 15808
rect 22784 15748 22788 15804
rect 22788 15748 22844 15804
rect 22844 15748 22848 15804
rect 22784 15744 22848 15748
rect 22864 15804 22928 15808
rect 22864 15748 22868 15804
rect 22868 15748 22924 15804
rect 22924 15748 22928 15804
rect 22864 15744 22928 15748
rect 37072 15804 37136 15808
rect 37072 15748 37076 15804
rect 37076 15748 37132 15804
rect 37132 15748 37136 15804
rect 37072 15744 37136 15748
rect 37152 15804 37216 15808
rect 37152 15748 37156 15804
rect 37156 15748 37212 15804
rect 37212 15748 37216 15804
rect 37152 15744 37216 15748
rect 37232 15804 37296 15808
rect 37232 15748 37236 15804
rect 37236 15748 37292 15804
rect 37292 15748 37296 15804
rect 37232 15744 37296 15748
rect 37312 15804 37376 15808
rect 37312 15748 37316 15804
rect 37316 15748 37372 15804
rect 37372 15748 37376 15804
rect 37312 15744 37376 15748
rect 51520 15804 51584 15808
rect 51520 15748 51524 15804
rect 51524 15748 51580 15804
rect 51580 15748 51584 15804
rect 51520 15744 51584 15748
rect 51600 15804 51664 15808
rect 51600 15748 51604 15804
rect 51604 15748 51660 15804
rect 51660 15748 51664 15804
rect 51600 15744 51664 15748
rect 51680 15804 51744 15808
rect 51680 15748 51684 15804
rect 51684 15748 51740 15804
rect 51740 15748 51744 15804
rect 51680 15744 51744 15748
rect 51760 15804 51824 15808
rect 51760 15748 51764 15804
rect 51764 15748 51820 15804
rect 51820 15748 51824 15804
rect 51760 15744 51824 15748
rect 15400 15260 15464 15264
rect 15400 15204 15404 15260
rect 15404 15204 15460 15260
rect 15460 15204 15464 15260
rect 15400 15200 15464 15204
rect 15480 15260 15544 15264
rect 15480 15204 15484 15260
rect 15484 15204 15540 15260
rect 15540 15204 15544 15260
rect 15480 15200 15544 15204
rect 15560 15260 15624 15264
rect 15560 15204 15564 15260
rect 15564 15204 15620 15260
rect 15620 15204 15624 15260
rect 15560 15200 15624 15204
rect 15640 15260 15704 15264
rect 15640 15204 15644 15260
rect 15644 15204 15700 15260
rect 15700 15204 15704 15260
rect 15640 15200 15704 15204
rect 29848 15260 29912 15264
rect 29848 15204 29852 15260
rect 29852 15204 29908 15260
rect 29908 15204 29912 15260
rect 29848 15200 29912 15204
rect 29928 15260 29992 15264
rect 29928 15204 29932 15260
rect 29932 15204 29988 15260
rect 29988 15204 29992 15260
rect 29928 15200 29992 15204
rect 30008 15260 30072 15264
rect 30008 15204 30012 15260
rect 30012 15204 30068 15260
rect 30068 15204 30072 15260
rect 30008 15200 30072 15204
rect 30088 15260 30152 15264
rect 30088 15204 30092 15260
rect 30092 15204 30148 15260
rect 30148 15204 30152 15260
rect 30088 15200 30152 15204
rect 44296 15260 44360 15264
rect 44296 15204 44300 15260
rect 44300 15204 44356 15260
rect 44356 15204 44360 15260
rect 44296 15200 44360 15204
rect 44376 15260 44440 15264
rect 44376 15204 44380 15260
rect 44380 15204 44436 15260
rect 44436 15204 44440 15260
rect 44376 15200 44440 15204
rect 44456 15260 44520 15264
rect 44456 15204 44460 15260
rect 44460 15204 44516 15260
rect 44516 15204 44520 15260
rect 44456 15200 44520 15204
rect 44536 15260 44600 15264
rect 44536 15204 44540 15260
rect 44540 15204 44596 15260
rect 44596 15204 44600 15260
rect 44536 15200 44600 15204
rect 8176 14716 8240 14720
rect 8176 14660 8180 14716
rect 8180 14660 8236 14716
rect 8236 14660 8240 14716
rect 8176 14656 8240 14660
rect 8256 14716 8320 14720
rect 8256 14660 8260 14716
rect 8260 14660 8316 14716
rect 8316 14660 8320 14716
rect 8256 14656 8320 14660
rect 8336 14716 8400 14720
rect 8336 14660 8340 14716
rect 8340 14660 8396 14716
rect 8396 14660 8400 14716
rect 8336 14656 8400 14660
rect 8416 14716 8480 14720
rect 8416 14660 8420 14716
rect 8420 14660 8476 14716
rect 8476 14660 8480 14716
rect 8416 14656 8480 14660
rect 22624 14716 22688 14720
rect 22624 14660 22628 14716
rect 22628 14660 22684 14716
rect 22684 14660 22688 14716
rect 22624 14656 22688 14660
rect 22704 14716 22768 14720
rect 22704 14660 22708 14716
rect 22708 14660 22764 14716
rect 22764 14660 22768 14716
rect 22704 14656 22768 14660
rect 22784 14716 22848 14720
rect 22784 14660 22788 14716
rect 22788 14660 22844 14716
rect 22844 14660 22848 14716
rect 22784 14656 22848 14660
rect 22864 14716 22928 14720
rect 22864 14660 22868 14716
rect 22868 14660 22924 14716
rect 22924 14660 22928 14716
rect 22864 14656 22928 14660
rect 37072 14716 37136 14720
rect 37072 14660 37076 14716
rect 37076 14660 37132 14716
rect 37132 14660 37136 14716
rect 37072 14656 37136 14660
rect 37152 14716 37216 14720
rect 37152 14660 37156 14716
rect 37156 14660 37212 14716
rect 37212 14660 37216 14716
rect 37152 14656 37216 14660
rect 37232 14716 37296 14720
rect 37232 14660 37236 14716
rect 37236 14660 37292 14716
rect 37292 14660 37296 14716
rect 37232 14656 37296 14660
rect 37312 14716 37376 14720
rect 37312 14660 37316 14716
rect 37316 14660 37372 14716
rect 37372 14660 37376 14716
rect 37312 14656 37376 14660
rect 51520 14716 51584 14720
rect 51520 14660 51524 14716
rect 51524 14660 51580 14716
rect 51580 14660 51584 14716
rect 51520 14656 51584 14660
rect 51600 14716 51664 14720
rect 51600 14660 51604 14716
rect 51604 14660 51660 14716
rect 51660 14660 51664 14716
rect 51600 14656 51664 14660
rect 51680 14716 51744 14720
rect 51680 14660 51684 14716
rect 51684 14660 51740 14716
rect 51740 14660 51744 14716
rect 51680 14656 51744 14660
rect 51760 14716 51824 14720
rect 51760 14660 51764 14716
rect 51764 14660 51820 14716
rect 51820 14660 51824 14716
rect 51760 14656 51824 14660
rect 15400 14172 15464 14176
rect 15400 14116 15404 14172
rect 15404 14116 15460 14172
rect 15460 14116 15464 14172
rect 15400 14112 15464 14116
rect 15480 14172 15544 14176
rect 15480 14116 15484 14172
rect 15484 14116 15540 14172
rect 15540 14116 15544 14172
rect 15480 14112 15544 14116
rect 15560 14172 15624 14176
rect 15560 14116 15564 14172
rect 15564 14116 15620 14172
rect 15620 14116 15624 14172
rect 15560 14112 15624 14116
rect 15640 14172 15704 14176
rect 15640 14116 15644 14172
rect 15644 14116 15700 14172
rect 15700 14116 15704 14172
rect 15640 14112 15704 14116
rect 29848 14172 29912 14176
rect 29848 14116 29852 14172
rect 29852 14116 29908 14172
rect 29908 14116 29912 14172
rect 29848 14112 29912 14116
rect 29928 14172 29992 14176
rect 29928 14116 29932 14172
rect 29932 14116 29988 14172
rect 29988 14116 29992 14172
rect 29928 14112 29992 14116
rect 30008 14172 30072 14176
rect 30008 14116 30012 14172
rect 30012 14116 30068 14172
rect 30068 14116 30072 14172
rect 30008 14112 30072 14116
rect 30088 14172 30152 14176
rect 30088 14116 30092 14172
rect 30092 14116 30148 14172
rect 30148 14116 30152 14172
rect 30088 14112 30152 14116
rect 44296 14172 44360 14176
rect 44296 14116 44300 14172
rect 44300 14116 44356 14172
rect 44356 14116 44360 14172
rect 44296 14112 44360 14116
rect 44376 14172 44440 14176
rect 44376 14116 44380 14172
rect 44380 14116 44436 14172
rect 44436 14116 44440 14172
rect 44376 14112 44440 14116
rect 44456 14172 44520 14176
rect 44456 14116 44460 14172
rect 44460 14116 44516 14172
rect 44516 14116 44520 14172
rect 44456 14112 44520 14116
rect 44536 14172 44600 14176
rect 44536 14116 44540 14172
rect 44540 14116 44596 14172
rect 44596 14116 44600 14172
rect 44536 14112 44600 14116
rect 8176 13628 8240 13632
rect 8176 13572 8180 13628
rect 8180 13572 8236 13628
rect 8236 13572 8240 13628
rect 8176 13568 8240 13572
rect 8256 13628 8320 13632
rect 8256 13572 8260 13628
rect 8260 13572 8316 13628
rect 8316 13572 8320 13628
rect 8256 13568 8320 13572
rect 8336 13628 8400 13632
rect 8336 13572 8340 13628
rect 8340 13572 8396 13628
rect 8396 13572 8400 13628
rect 8336 13568 8400 13572
rect 8416 13628 8480 13632
rect 8416 13572 8420 13628
rect 8420 13572 8476 13628
rect 8476 13572 8480 13628
rect 8416 13568 8480 13572
rect 22624 13628 22688 13632
rect 22624 13572 22628 13628
rect 22628 13572 22684 13628
rect 22684 13572 22688 13628
rect 22624 13568 22688 13572
rect 22704 13628 22768 13632
rect 22704 13572 22708 13628
rect 22708 13572 22764 13628
rect 22764 13572 22768 13628
rect 22704 13568 22768 13572
rect 22784 13628 22848 13632
rect 22784 13572 22788 13628
rect 22788 13572 22844 13628
rect 22844 13572 22848 13628
rect 22784 13568 22848 13572
rect 22864 13628 22928 13632
rect 22864 13572 22868 13628
rect 22868 13572 22924 13628
rect 22924 13572 22928 13628
rect 22864 13568 22928 13572
rect 37072 13628 37136 13632
rect 37072 13572 37076 13628
rect 37076 13572 37132 13628
rect 37132 13572 37136 13628
rect 37072 13568 37136 13572
rect 37152 13628 37216 13632
rect 37152 13572 37156 13628
rect 37156 13572 37212 13628
rect 37212 13572 37216 13628
rect 37152 13568 37216 13572
rect 37232 13628 37296 13632
rect 37232 13572 37236 13628
rect 37236 13572 37292 13628
rect 37292 13572 37296 13628
rect 37232 13568 37296 13572
rect 37312 13628 37376 13632
rect 37312 13572 37316 13628
rect 37316 13572 37372 13628
rect 37372 13572 37376 13628
rect 37312 13568 37376 13572
rect 51520 13628 51584 13632
rect 51520 13572 51524 13628
rect 51524 13572 51580 13628
rect 51580 13572 51584 13628
rect 51520 13568 51584 13572
rect 51600 13628 51664 13632
rect 51600 13572 51604 13628
rect 51604 13572 51660 13628
rect 51660 13572 51664 13628
rect 51600 13568 51664 13572
rect 51680 13628 51744 13632
rect 51680 13572 51684 13628
rect 51684 13572 51740 13628
rect 51740 13572 51744 13628
rect 51680 13568 51744 13572
rect 51760 13628 51824 13632
rect 51760 13572 51764 13628
rect 51764 13572 51820 13628
rect 51820 13572 51824 13628
rect 51760 13568 51824 13572
rect 15400 13084 15464 13088
rect 15400 13028 15404 13084
rect 15404 13028 15460 13084
rect 15460 13028 15464 13084
rect 15400 13024 15464 13028
rect 15480 13084 15544 13088
rect 15480 13028 15484 13084
rect 15484 13028 15540 13084
rect 15540 13028 15544 13084
rect 15480 13024 15544 13028
rect 15560 13084 15624 13088
rect 15560 13028 15564 13084
rect 15564 13028 15620 13084
rect 15620 13028 15624 13084
rect 15560 13024 15624 13028
rect 15640 13084 15704 13088
rect 15640 13028 15644 13084
rect 15644 13028 15700 13084
rect 15700 13028 15704 13084
rect 15640 13024 15704 13028
rect 29848 13084 29912 13088
rect 29848 13028 29852 13084
rect 29852 13028 29908 13084
rect 29908 13028 29912 13084
rect 29848 13024 29912 13028
rect 29928 13084 29992 13088
rect 29928 13028 29932 13084
rect 29932 13028 29988 13084
rect 29988 13028 29992 13084
rect 29928 13024 29992 13028
rect 30008 13084 30072 13088
rect 30008 13028 30012 13084
rect 30012 13028 30068 13084
rect 30068 13028 30072 13084
rect 30008 13024 30072 13028
rect 30088 13084 30152 13088
rect 30088 13028 30092 13084
rect 30092 13028 30148 13084
rect 30148 13028 30152 13084
rect 30088 13024 30152 13028
rect 44296 13084 44360 13088
rect 44296 13028 44300 13084
rect 44300 13028 44356 13084
rect 44356 13028 44360 13084
rect 44296 13024 44360 13028
rect 44376 13084 44440 13088
rect 44376 13028 44380 13084
rect 44380 13028 44436 13084
rect 44436 13028 44440 13084
rect 44376 13024 44440 13028
rect 44456 13084 44520 13088
rect 44456 13028 44460 13084
rect 44460 13028 44516 13084
rect 44516 13028 44520 13084
rect 44456 13024 44520 13028
rect 44536 13084 44600 13088
rect 44536 13028 44540 13084
rect 44540 13028 44596 13084
rect 44596 13028 44600 13084
rect 44536 13024 44600 13028
rect 8176 12540 8240 12544
rect 8176 12484 8180 12540
rect 8180 12484 8236 12540
rect 8236 12484 8240 12540
rect 8176 12480 8240 12484
rect 8256 12540 8320 12544
rect 8256 12484 8260 12540
rect 8260 12484 8316 12540
rect 8316 12484 8320 12540
rect 8256 12480 8320 12484
rect 8336 12540 8400 12544
rect 8336 12484 8340 12540
rect 8340 12484 8396 12540
rect 8396 12484 8400 12540
rect 8336 12480 8400 12484
rect 8416 12540 8480 12544
rect 8416 12484 8420 12540
rect 8420 12484 8476 12540
rect 8476 12484 8480 12540
rect 8416 12480 8480 12484
rect 22624 12540 22688 12544
rect 22624 12484 22628 12540
rect 22628 12484 22684 12540
rect 22684 12484 22688 12540
rect 22624 12480 22688 12484
rect 22704 12540 22768 12544
rect 22704 12484 22708 12540
rect 22708 12484 22764 12540
rect 22764 12484 22768 12540
rect 22704 12480 22768 12484
rect 22784 12540 22848 12544
rect 22784 12484 22788 12540
rect 22788 12484 22844 12540
rect 22844 12484 22848 12540
rect 22784 12480 22848 12484
rect 22864 12540 22928 12544
rect 22864 12484 22868 12540
rect 22868 12484 22924 12540
rect 22924 12484 22928 12540
rect 22864 12480 22928 12484
rect 37072 12540 37136 12544
rect 37072 12484 37076 12540
rect 37076 12484 37132 12540
rect 37132 12484 37136 12540
rect 37072 12480 37136 12484
rect 37152 12540 37216 12544
rect 37152 12484 37156 12540
rect 37156 12484 37212 12540
rect 37212 12484 37216 12540
rect 37152 12480 37216 12484
rect 37232 12540 37296 12544
rect 37232 12484 37236 12540
rect 37236 12484 37292 12540
rect 37292 12484 37296 12540
rect 37232 12480 37296 12484
rect 37312 12540 37376 12544
rect 37312 12484 37316 12540
rect 37316 12484 37372 12540
rect 37372 12484 37376 12540
rect 37312 12480 37376 12484
rect 51520 12540 51584 12544
rect 51520 12484 51524 12540
rect 51524 12484 51580 12540
rect 51580 12484 51584 12540
rect 51520 12480 51584 12484
rect 51600 12540 51664 12544
rect 51600 12484 51604 12540
rect 51604 12484 51660 12540
rect 51660 12484 51664 12540
rect 51600 12480 51664 12484
rect 51680 12540 51744 12544
rect 51680 12484 51684 12540
rect 51684 12484 51740 12540
rect 51740 12484 51744 12540
rect 51680 12480 51744 12484
rect 51760 12540 51824 12544
rect 51760 12484 51764 12540
rect 51764 12484 51820 12540
rect 51820 12484 51824 12540
rect 51760 12480 51824 12484
rect 15400 11996 15464 12000
rect 15400 11940 15404 11996
rect 15404 11940 15460 11996
rect 15460 11940 15464 11996
rect 15400 11936 15464 11940
rect 15480 11996 15544 12000
rect 15480 11940 15484 11996
rect 15484 11940 15540 11996
rect 15540 11940 15544 11996
rect 15480 11936 15544 11940
rect 15560 11996 15624 12000
rect 15560 11940 15564 11996
rect 15564 11940 15620 11996
rect 15620 11940 15624 11996
rect 15560 11936 15624 11940
rect 15640 11996 15704 12000
rect 15640 11940 15644 11996
rect 15644 11940 15700 11996
rect 15700 11940 15704 11996
rect 15640 11936 15704 11940
rect 29848 11996 29912 12000
rect 29848 11940 29852 11996
rect 29852 11940 29908 11996
rect 29908 11940 29912 11996
rect 29848 11936 29912 11940
rect 29928 11996 29992 12000
rect 29928 11940 29932 11996
rect 29932 11940 29988 11996
rect 29988 11940 29992 11996
rect 29928 11936 29992 11940
rect 30008 11996 30072 12000
rect 30008 11940 30012 11996
rect 30012 11940 30068 11996
rect 30068 11940 30072 11996
rect 30008 11936 30072 11940
rect 30088 11996 30152 12000
rect 30088 11940 30092 11996
rect 30092 11940 30148 11996
rect 30148 11940 30152 11996
rect 30088 11936 30152 11940
rect 44296 11996 44360 12000
rect 44296 11940 44300 11996
rect 44300 11940 44356 11996
rect 44356 11940 44360 11996
rect 44296 11936 44360 11940
rect 44376 11996 44440 12000
rect 44376 11940 44380 11996
rect 44380 11940 44436 11996
rect 44436 11940 44440 11996
rect 44376 11936 44440 11940
rect 44456 11996 44520 12000
rect 44456 11940 44460 11996
rect 44460 11940 44516 11996
rect 44516 11940 44520 11996
rect 44456 11936 44520 11940
rect 44536 11996 44600 12000
rect 44536 11940 44540 11996
rect 44540 11940 44596 11996
rect 44596 11940 44600 11996
rect 44536 11936 44600 11940
rect 8176 11452 8240 11456
rect 8176 11396 8180 11452
rect 8180 11396 8236 11452
rect 8236 11396 8240 11452
rect 8176 11392 8240 11396
rect 8256 11452 8320 11456
rect 8256 11396 8260 11452
rect 8260 11396 8316 11452
rect 8316 11396 8320 11452
rect 8256 11392 8320 11396
rect 8336 11452 8400 11456
rect 8336 11396 8340 11452
rect 8340 11396 8396 11452
rect 8396 11396 8400 11452
rect 8336 11392 8400 11396
rect 8416 11452 8480 11456
rect 8416 11396 8420 11452
rect 8420 11396 8476 11452
rect 8476 11396 8480 11452
rect 8416 11392 8480 11396
rect 22624 11452 22688 11456
rect 22624 11396 22628 11452
rect 22628 11396 22684 11452
rect 22684 11396 22688 11452
rect 22624 11392 22688 11396
rect 22704 11452 22768 11456
rect 22704 11396 22708 11452
rect 22708 11396 22764 11452
rect 22764 11396 22768 11452
rect 22704 11392 22768 11396
rect 22784 11452 22848 11456
rect 22784 11396 22788 11452
rect 22788 11396 22844 11452
rect 22844 11396 22848 11452
rect 22784 11392 22848 11396
rect 22864 11452 22928 11456
rect 22864 11396 22868 11452
rect 22868 11396 22924 11452
rect 22924 11396 22928 11452
rect 22864 11392 22928 11396
rect 37072 11452 37136 11456
rect 37072 11396 37076 11452
rect 37076 11396 37132 11452
rect 37132 11396 37136 11452
rect 37072 11392 37136 11396
rect 37152 11452 37216 11456
rect 37152 11396 37156 11452
rect 37156 11396 37212 11452
rect 37212 11396 37216 11452
rect 37152 11392 37216 11396
rect 37232 11452 37296 11456
rect 37232 11396 37236 11452
rect 37236 11396 37292 11452
rect 37292 11396 37296 11452
rect 37232 11392 37296 11396
rect 37312 11452 37376 11456
rect 37312 11396 37316 11452
rect 37316 11396 37372 11452
rect 37372 11396 37376 11452
rect 37312 11392 37376 11396
rect 51520 11452 51584 11456
rect 51520 11396 51524 11452
rect 51524 11396 51580 11452
rect 51580 11396 51584 11452
rect 51520 11392 51584 11396
rect 51600 11452 51664 11456
rect 51600 11396 51604 11452
rect 51604 11396 51660 11452
rect 51660 11396 51664 11452
rect 51600 11392 51664 11396
rect 51680 11452 51744 11456
rect 51680 11396 51684 11452
rect 51684 11396 51740 11452
rect 51740 11396 51744 11452
rect 51680 11392 51744 11396
rect 51760 11452 51824 11456
rect 51760 11396 51764 11452
rect 51764 11396 51820 11452
rect 51820 11396 51824 11452
rect 51760 11392 51824 11396
rect 15400 10908 15464 10912
rect 15400 10852 15404 10908
rect 15404 10852 15460 10908
rect 15460 10852 15464 10908
rect 15400 10848 15464 10852
rect 15480 10908 15544 10912
rect 15480 10852 15484 10908
rect 15484 10852 15540 10908
rect 15540 10852 15544 10908
rect 15480 10848 15544 10852
rect 15560 10908 15624 10912
rect 15560 10852 15564 10908
rect 15564 10852 15620 10908
rect 15620 10852 15624 10908
rect 15560 10848 15624 10852
rect 15640 10908 15704 10912
rect 15640 10852 15644 10908
rect 15644 10852 15700 10908
rect 15700 10852 15704 10908
rect 15640 10848 15704 10852
rect 29848 10908 29912 10912
rect 29848 10852 29852 10908
rect 29852 10852 29908 10908
rect 29908 10852 29912 10908
rect 29848 10848 29912 10852
rect 29928 10908 29992 10912
rect 29928 10852 29932 10908
rect 29932 10852 29988 10908
rect 29988 10852 29992 10908
rect 29928 10848 29992 10852
rect 30008 10908 30072 10912
rect 30008 10852 30012 10908
rect 30012 10852 30068 10908
rect 30068 10852 30072 10908
rect 30008 10848 30072 10852
rect 30088 10908 30152 10912
rect 30088 10852 30092 10908
rect 30092 10852 30148 10908
rect 30148 10852 30152 10908
rect 30088 10848 30152 10852
rect 44296 10908 44360 10912
rect 44296 10852 44300 10908
rect 44300 10852 44356 10908
rect 44356 10852 44360 10908
rect 44296 10848 44360 10852
rect 44376 10908 44440 10912
rect 44376 10852 44380 10908
rect 44380 10852 44436 10908
rect 44436 10852 44440 10908
rect 44376 10848 44440 10852
rect 44456 10908 44520 10912
rect 44456 10852 44460 10908
rect 44460 10852 44516 10908
rect 44516 10852 44520 10908
rect 44456 10848 44520 10852
rect 44536 10908 44600 10912
rect 44536 10852 44540 10908
rect 44540 10852 44596 10908
rect 44596 10852 44600 10908
rect 44536 10848 44600 10852
rect 8176 10364 8240 10368
rect 8176 10308 8180 10364
rect 8180 10308 8236 10364
rect 8236 10308 8240 10364
rect 8176 10304 8240 10308
rect 8256 10364 8320 10368
rect 8256 10308 8260 10364
rect 8260 10308 8316 10364
rect 8316 10308 8320 10364
rect 8256 10304 8320 10308
rect 8336 10364 8400 10368
rect 8336 10308 8340 10364
rect 8340 10308 8396 10364
rect 8396 10308 8400 10364
rect 8336 10304 8400 10308
rect 8416 10364 8480 10368
rect 8416 10308 8420 10364
rect 8420 10308 8476 10364
rect 8476 10308 8480 10364
rect 8416 10304 8480 10308
rect 22624 10364 22688 10368
rect 22624 10308 22628 10364
rect 22628 10308 22684 10364
rect 22684 10308 22688 10364
rect 22624 10304 22688 10308
rect 22704 10364 22768 10368
rect 22704 10308 22708 10364
rect 22708 10308 22764 10364
rect 22764 10308 22768 10364
rect 22704 10304 22768 10308
rect 22784 10364 22848 10368
rect 22784 10308 22788 10364
rect 22788 10308 22844 10364
rect 22844 10308 22848 10364
rect 22784 10304 22848 10308
rect 22864 10364 22928 10368
rect 22864 10308 22868 10364
rect 22868 10308 22924 10364
rect 22924 10308 22928 10364
rect 22864 10304 22928 10308
rect 37072 10364 37136 10368
rect 37072 10308 37076 10364
rect 37076 10308 37132 10364
rect 37132 10308 37136 10364
rect 37072 10304 37136 10308
rect 37152 10364 37216 10368
rect 37152 10308 37156 10364
rect 37156 10308 37212 10364
rect 37212 10308 37216 10364
rect 37152 10304 37216 10308
rect 37232 10364 37296 10368
rect 37232 10308 37236 10364
rect 37236 10308 37292 10364
rect 37292 10308 37296 10364
rect 37232 10304 37296 10308
rect 37312 10364 37376 10368
rect 37312 10308 37316 10364
rect 37316 10308 37372 10364
rect 37372 10308 37376 10364
rect 37312 10304 37376 10308
rect 51520 10364 51584 10368
rect 51520 10308 51524 10364
rect 51524 10308 51580 10364
rect 51580 10308 51584 10364
rect 51520 10304 51584 10308
rect 51600 10364 51664 10368
rect 51600 10308 51604 10364
rect 51604 10308 51660 10364
rect 51660 10308 51664 10364
rect 51600 10304 51664 10308
rect 51680 10364 51744 10368
rect 51680 10308 51684 10364
rect 51684 10308 51740 10364
rect 51740 10308 51744 10364
rect 51680 10304 51744 10308
rect 51760 10364 51824 10368
rect 51760 10308 51764 10364
rect 51764 10308 51820 10364
rect 51820 10308 51824 10364
rect 51760 10304 51824 10308
rect 15400 9820 15464 9824
rect 15400 9764 15404 9820
rect 15404 9764 15460 9820
rect 15460 9764 15464 9820
rect 15400 9760 15464 9764
rect 15480 9820 15544 9824
rect 15480 9764 15484 9820
rect 15484 9764 15540 9820
rect 15540 9764 15544 9820
rect 15480 9760 15544 9764
rect 15560 9820 15624 9824
rect 15560 9764 15564 9820
rect 15564 9764 15620 9820
rect 15620 9764 15624 9820
rect 15560 9760 15624 9764
rect 15640 9820 15704 9824
rect 15640 9764 15644 9820
rect 15644 9764 15700 9820
rect 15700 9764 15704 9820
rect 15640 9760 15704 9764
rect 29848 9820 29912 9824
rect 29848 9764 29852 9820
rect 29852 9764 29908 9820
rect 29908 9764 29912 9820
rect 29848 9760 29912 9764
rect 29928 9820 29992 9824
rect 29928 9764 29932 9820
rect 29932 9764 29988 9820
rect 29988 9764 29992 9820
rect 29928 9760 29992 9764
rect 30008 9820 30072 9824
rect 30008 9764 30012 9820
rect 30012 9764 30068 9820
rect 30068 9764 30072 9820
rect 30008 9760 30072 9764
rect 30088 9820 30152 9824
rect 30088 9764 30092 9820
rect 30092 9764 30148 9820
rect 30148 9764 30152 9820
rect 30088 9760 30152 9764
rect 44296 9820 44360 9824
rect 44296 9764 44300 9820
rect 44300 9764 44356 9820
rect 44356 9764 44360 9820
rect 44296 9760 44360 9764
rect 44376 9820 44440 9824
rect 44376 9764 44380 9820
rect 44380 9764 44436 9820
rect 44436 9764 44440 9820
rect 44376 9760 44440 9764
rect 44456 9820 44520 9824
rect 44456 9764 44460 9820
rect 44460 9764 44516 9820
rect 44516 9764 44520 9820
rect 44456 9760 44520 9764
rect 44536 9820 44600 9824
rect 44536 9764 44540 9820
rect 44540 9764 44596 9820
rect 44596 9764 44600 9820
rect 44536 9760 44600 9764
rect 8176 9276 8240 9280
rect 8176 9220 8180 9276
rect 8180 9220 8236 9276
rect 8236 9220 8240 9276
rect 8176 9216 8240 9220
rect 8256 9276 8320 9280
rect 8256 9220 8260 9276
rect 8260 9220 8316 9276
rect 8316 9220 8320 9276
rect 8256 9216 8320 9220
rect 8336 9276 8400 9280
rect 8336 9220 8340 9276
rect 8340 9220 8396 9276
rect 8396 9220 8400 9276
rect 8336 9216 8400 9220
rect 8416 9276 8480 9280
rect 8416 9220 8420 9276
rect 8420 9220 8476 9276
rect 8476 9220 8480 9276
rect 8416 9216 8480 9220
rect 22624 9276 22688 9280
rect 22624 9220 22628 9276
rect 22628 9220 22684 9276
rect 22684 9220 22688 9276
rect 22624 9216 22688 9220
rect 22704 9276 22768 9280
rect 22704 9220 22708 9276
rect 22708 9220 22764 9276
rect 22764 9220 22768 9276
rect 22704 9216 22768 9220
rect 22784 9276 22848 9280
rect 22784 9220 22788 9276
rect 22788 9220 22844 9276
rect 22844 9220 22848 9276
rect 22784 9216 22848 9220
rect 22864 9276 22928 9280
rect 22864 9220 22868 9276
rect 22868 9220 22924 9276
rect 22924 9220 22928 9276
rect 22864 9216 22928 9220
rect 37072 9276 37136 9280
rect 37072 9220 37076 9276
rect 37076 9220 37132 9276
rect 37132 9220 37136 9276
rect 37072 9216 37136 9220
rect 37152 9276 37216 9280
rect 37152 9220 37156 9276
rect 37156 9220 37212 9276
rect 37212 9220 37216 9276
rect 37152 9216 37216 9220
rect 37232 9276 37296 9280
rect 37232 9220 37236 9276
rect 37236 9220 37292 9276
rect 37292 9220 37296 9276
rect 37232 9216 37296 9220
rect 37312 9276 37376 9280
rect 37312 9220 37316 9276
rect 37316 9220 37372 9276
rect 37372 9220 37376 9276
rect 37312 9216 37376 9220
rect 51520 9276 51584 9280
rect 51520 9220 51524 9276
rect 51524 9220 51580 9276
rect 51580 9220 51584 9276
rect 51520 9216 51584 9220
rect 51600 9276 51664 9280
rect 51600 9220 51604 9276
rect 51604 9220 51660 9276
rect 51660 9220 51664 9276
rect 51600 9216 51664 9220
rect 51680 9276 51744 9280
rect 51680 9220 51684 9276
rect 51684 9220 51740 9276
rect 51740 9220 51744 9276
rect 51680 9216 51744 9220
rect 51760 9276 51824 9280
rect 51760 9220 51764 9276
rect 51764 9220 51820 9276
rect 51820 9220 51824 9276
rect 51760 9216 51824 9220
rect 15400 8732 15464 8736
rect 15400 8676 15404 8732
rect 15404 8676 15460 8732
rect 15460 8676 15464 8732
rect 15400 8672 15464 8676
rect 15480 8732 15544 8736
rect 15480 8676 15484 8732
rect 15484 8676 15540 8732
rect 15540 8676 15544 8732
rect 15480 8672 15544 8676
rect 15560 8732 15624 8736
rect 15560 8676 15564 8732
rect 15564 8676 15620 8732
rect 15620 8676 15624 8732
rect 15560 8672 15624 8676
rect 15640 8732 15704 8736
rect 15640 8676 15644 8732
rect 15644 8676 15700 8732
rect 15700 8676 15704 8732
rect 15640 8672 15704 8676
rect 29848 8732 29912 8736
rect 29848 8676 29852 8732
rect 29852 8676 29908 8732
rect 29908 8676 29912 8732
rect 29848 8672 29912 8676
rect 29928 8732 29992 8736
rect 29928 8676 29932 8732
rect 29932 8676 29988 8732
rect 29988 8676 29992 8732
rect 29928 8672 29992 8676
rect 30008 8732 30072 8736
rect 30008 8676 30012 8732
rect 30012 8676 30068 8732
rect 30068 8676 30072 8732
rect 30008 8672 30072 8676
rect 30088 8732 30152 8736
rect 30088 8676 30092 8732
rect 30092 8676 30148 8732
rect 30148 8676 30152 8732
rect 30088 8672 30152 8676
rect 44296 8732 44360 8736
rect 44296 8676 44300 8732
rect 44300 8676 44356 8732
rect 44356 8676 44360 8732
rect 44296 8672 44360 8676
rect 44376 8732 44440 8736
rect 44376 8676 44380 8732
rect 44380 8676 44436 8732
rect 44436 8676 44440 8732
rect 44376 8672 44440 8676
rect 44456 8732 44520 8736
rect 44456 8676 44460 8732
rect 44460 8676 44516 8732
rect 44516 8676 44520 8732
rect 44456 8672 44520 8676
rect 44536 8732 44600 8736
rect 44536 8676 44540 8732
rect 44540 8676 44596 8732
rect 44596 8676 44600 8732
rect 44536 8672 44600 8676
rect 8176 8188 8240 8192
rect 8176 8132 8180 8188
rect 8180 8132 8236 8188
rect 8236 8132 8240 8188
rect 8176 8128 8240 8132
rect 8256 8188 8320 8192
rect 8256 8132 8260 8188
rect 8260 8132 8316 8188
rect 8316 8132 8320 8188
rect 8256 8128 8320 8132
rect 8336 8188 8400 8192
rect 8336 8132 8340 8188
rect 8340 8132 8396 8188
rect 8396 8132 8400 8188
rect 8336 8128 8400 8132
rect 8416 8188 8480 8192
rect 8416 8132 8420 8188
rect 8420 8132 8476 8188
rect 8476 8132 8480 8188
rect 8416 8128 8480 8132
rect 22624 8188 22688 8192
rect 22624 8132 22628 8188
rect 22628 8132 22684 8188
rect 22684 8132 22688 8188
rect 22624 8128 22688 8132
rect 22704 8188 22768 8192
rect 22704 8132 22708 8188
rect 22708 8132 22764 8188
rect 22764 8132 22768 8188
rect 22704 8128 22768 8132
rect 22784 8188 22848 8192
rect 22784 8132 22788 8188
rect 22788 8132 22844 8188
rect 22844 8132 22848 8188
rect 22784 8128 22848 8132
rect 22864 8188 22928 8192
rect 22864 8132 22868 8188
rect 22868 8132 22924 8188
rect 22924 8132 22928 8188
rect 22864 8128 22928 8132
rect 37072 8188 37136 8192
rect 37072 8132 37076 8188
rect 37076 8132 37132 8188
rect 37132 8132 37136 8188
rect 37072 8128 37136 8132
rect 37152 8188 37216 8192
rect 37152 8132 37156 8188
rect 37156 8132 37212 8188
rect 37212 8132 37216 8188
rect 37152 8128 37216 8132
rect 37232 8188 37296 8192
rect 37232 8132 37236 8188
rect 37236 8132 37292 8188
rect 37292 8132 37296 8188
rect 37232 8128 37296 8132
rect 37312 8188 37376 8192
rect 37312 8132 37316 8188
rect 37316 8132 37372 8188
rect 37372 8132 37376 8188
rect 37312 8128 37376 8132
rect 51520 8188 51584 8192
rect 51520 8132 51524 8188
rect 51524 8132 51580 8188
rect 51580 8132 51584 8188
rect 51520 8128 51584 8132
rect 51600 8188 51664 8192
rect 51600 8132 51604 8188
rect 51604 8132 51660 8188
rect 51660 8132 51664 8188
rect 51600 8128 51664 8132
rect 51680 8188 51744 8192
rect 51680 8132 51684 8188
rect 51684 8132 51740 8188
rect 51740 8132 51744 8188
rect 51680 8128 51744 8132
rect 51760 8188 51824 8192
rect 51760 8132 51764 8188
rect 51764 8132 51820 8188
rect 51820 8132 51824 8188
rect 51760 8128 51824 8132
rect 15400 7644 15464 7648
rect 15400 7588 15404 7644
rect 15404 7588 15460 7644
rect 15460 7588 15464 7644
rect 15400 7584 15464 7588
rect 15480 7644 15544 7648
rect 15480 7588 15484 7644
rect 15484 7588 15540 7644
rect 15540 7588 15544 7644
rect 15480 7584 15544 7588
rect 15560 7644 15624 7648
rect 15560 7588 15564 7644
rect 15564 7588 15620 7644
rect 15620 7588 15624 7644
rect 15560 7584 15624 7588
rect 15640 7644 15704 7648
rect 15640 7588 15644 7644
rect 15644 7588 15700 7644
rect 15700 7588 15704 7644
rect 15640 7584 15704 7588
rect 29848 7644 29912 7648
rect 29848 7588 29852 7644
rect 29852 7588 29908 7644
rect 29908 7588 29912 7644
rect 29848 7584 29912 7588
rect 29928 7644 29992 7648
rect 29928 7588 29932 7644
rect 29932 7588 29988 7644
rect 29988 7588 29992 7644
rect 29928 7584 29992 7588
rect 30008 7644 30072 7648
rect 30008 7588 30012 7644
rect 30012 7588 30068 7644
rect 30068 7588 30072 7644
rect 30008 7584 30072 7588
rect 30088 7644 30152 7648
rect 30088 7588 30092 7644
rect 30092 7588 30148 7644
rect 30148 7588 30152 7644
rect 30088 7584 30152 7588
rect 44296 7644 44360 7648
rect 44296 7588 44300 7644
rect 44300 7588 44356 7644
rect 44356 7588 44360 7644
rect 44296 7584 44360 7588
rect 44376 7644 44440 7648
rect 44376 7588 44380 7644
rect 44380 7588 44436 7644
rect 44436 7588 44440 7644
rect 44376 7584 44440 7588
rect 44456 7644 44520 7648
rect 44456 7588 44460 7644
rect 44460 7588 44516 7644
rect 44516 7588 44520 7644
rect 44456 7584 44520 7588
rect 44536 7644 44600 7648
rect 44536 7588 44540 7644
rect 44540 7588 44596 7644
rect 44596 7588 44600 7644
rect 44536 7584 44600 7588
rect 8176 7100 8240 7104
rect 8176 7044 8180 7100
rect 8180 7044 8236 7100
rect 8236 7044 8240 7100
rect 8176 7040 8240 7044
rect 8256 7100 8320 7104
rect 8256 7044 8260 7100
rect 8260 7044 8316 7100
rect 8316 7044 8320 7100
rect 8256 7040 8320 7044
rect 8336 7100 8400 7104
rect 8336 7044 8340 7100
rect 8340 7044 8396 7100
rect 8396 7044 8400 7100
rect 8336 7040 8400 7044
rect 8416 7100 8480 7104
rect 8416 7044 8420 7100
rect 8420 7044 8476 7100
rect 8476 7044 8480 7100
rect 8416 7040 8480 7044
rect 22624 7100 22688 7104
rect 22624 7044 22628 7100
rect 22628 7044 22684 7100
rect 22684 7044 22688 7100
rect 22624 7040 22688 7044
rect 22704 7100 22768 7104
rect 22704 7044 22708 7100
rect 22708 7044 22764 7100
rect 22764 7044 22768 7100
rect 22704 7040 22768 7044
rect 22784 7100 22848 7104
rect 22784 7044 22788 7100
rect 22788 7044 22844 7100
rect 22844 7044 22848 7100
rect 22784 7040 22848 7044
rect 22864 7100 22928 7104
rect 22864 7044 22868 7100
rect 22868 7044 22924 7100
rect 22924 7044 22928 7100
rect 22864 7040 22928 7044
rect 37072 7100 37136 7104
rect 37072 7044 37076 7100
rect 37076 7044 37132 7100
rect 37132 7044 37136 7100
rect 37072 7040 37136 7044
rect 37152 7100 37216 7104
rect 37152 7044 37156 7100
rect 37156 7044 37212 7100
rect 37212 7044 37216 7100
rect 37152 7040 37216 7044
rect 37232 7100 37296 7104
rect 37232 7044 37236 7100
rect 37236 7044 37292 7100
rect 37292 7044 37296 7100
rect 37232 7040 37296 7044
rect 37312 7100 37376 7104
rect 37312 7044 37316 7100
rect 37316 7044 37372 7100
rect 37372 7044 37376 7100
rect 37312 7040 37376 7044
rect 51520 7100 51584 7104
rect 51520 7044 51524 7100
rect 51524 7044 51580 7100
rect 51580 7044 51584 7100
rect 51520 7040 51584 7044
rect 51600 7100 51664 7104
rect 51600 7044 51604 7100
rect 51604 7044 51660 7100
rect 51660 7044 51664 7100
rect 51600 7040 51664 7044
rect 51680 7100 51744 7104
rect 51680 7044 51684 7100
rect 51684 7044 51740 7100
rect 51740 7044 51744 7100
rect 51680 7040 51744 7044
rect 51760 7100 51824 7104
rect 51760 7044 51764 7100
rect 51764 7044 51820 7100
rect 51820 7044 51824 7100
rect 51760 7040 51824 7044
rect 15400 6556 15464 6560
rect 15400 6500 15404 6556
rect 15404 6500 15460 6556
rect 15460 6500 15464 6556
rect 15400 6496 15464 6500
rect 15480 6556 15544 6560
rect 15480 6500 15484 6556
rect 15484 6500 15540 6556
rect 15540 6500 15544 6556
rect 15480 6496 15544 6500
rect 15560 6556 15624 6560
rect 15560 6500 15564 6556
rect 15564 6500 15620 6556
rect 15620 6500 15624 6556
rect 15560 6496 15624 6500
rect 15640 6556 15704 6560
rect 15640 6500 15644 6556
rect 15644 6500 15700 6556
rect 15700 6500 15704 6556
rect 15640 6496 15704 6500
rect 29848 6556 29912 6560
rect 29848 6500 29852 6556
rect 29852 6500 29908 6556
rect 29908 6500 29912 6556
rect 29848 6496 29912 6500
rect 29928 6556 29992 6560
rect 29928 6500 29932 6556
rect 29932 6500 29988 6556
rect 29988 6500 29992 6556
rect 29928 6496 29992 6500
rect 30008 6556 30072 6560
rect 30008 6500 30012 6556
rect 30012 6500 30068 6556
rect 30068 6500 30072 6556
rect 30008 6496 30072 6500
rect 30088 6556 30152 6560
rect 30088 6500 30092 6556
rect 30092 6500 30148 6556
rect 30148 6500 30152 6556
rect 30088 6496 30152 6500
rect 44296 6556 44360 6560
rect 44296 6500 44300 6556
rect 44300 6500 44356 6556
rect 44356 6500 44360 6556
rect 44296 6496 44360 6500
rect 44376 6556 44440 6560
rect 44376 6500 44380 6556
rect 44380 6500 44436 6556
rect 44436 6500 44440 6556
rect 44376 6496 44440 6500
rect 44456 6556 44520 6560
rect 44456 6500 44460 6556
rect 44460 6500 44516 6556
rect 44516 6500 44520 6556
rect 44456 6496 44520 6500
rect 44536 6556 44600 6560
rect 44536 6500 44540 6556
rect 44540 6500 44596 6556
rect 44596 6500 44600 6556
rect 44536 6496 44600 6500
rect 8176 6012 8240 6016
rect 8176 5956 8180 6012
rect 8180 5956 8236 6012
rect 8236 5956 8240 6012
rect 8176 5952 8240 5956
rect 8256 6012 8320 6016
rect 8256 5956 8260 6012
rect 8260 5956 8316 6012
rect 8316 5956 8320 6012
rect 8256 5952 8320 5956
rect 8336 6012 8400 6016
rect 8336 5956 8340 6012
rect 8340 5956 8396 6012
rect 8396 5956 8400 6012
rect 8336 5952 8400 5956
rect 8416 6012 8480 6016
rect 8416 5956 8420 6012
rect 8420 5956 8476 6012
rect 8476 5956 8480 6012
rect 8416 5952 8480 5956
rect 22624 6012 22688 6016
rect 22624 5956 22628 6012
rect 22628 5956 22684 6012
rect 22684 5956 22688 6012
rect 22624 5952 22688 5956
rect 22704 6012 22768 6016
rect 22704 5956 22708 6012
rect 22708 5956 22764 6012
rect 22764 5956 22768 6012
rect 22704 5952 22768 5956
rect 22784 6012 22848 6016
rect 22784 5956 22788 6012
rect 22788 5956 22844 6012
rect 22844 5956 22848 6012
rect 22784 5952 22848 5956
rect 22864 6012 22928 6016
rect 22864 5956 22868 6012
rect 22868 5956 22924 6012
rect 22924 5956 22928 6012
rect 22864 5952 22928 5956
rect 37072 6012 37136 6016
rect 37072 5956 37076 6012
rect 37076 5956 37132 6012
rect 37132 5956 37136 6012
rect 37072 5952 37136 5956
rect 37152 6012 37216 6016
rect 37152 5956 37156 6012
rect 37156 5956 37212 6012
rect 37212 5956 37216 6012
rect 37152 5952 37216 5956
rect 37232 6012 37296 6016
rect 37232 5956 37236 6012
rect 37236 5956 37292 6012
rect 37292 5956 37296 6012
rect 37232 5952 37296 5956
rect 37312 6012 37376 6016
rect 37312 5956 37316 6012
rect 37316 5956 37372 6012
rect 37372 5956 37376 6012
rect 37312 5952 37376 5956
rect 51520 6012 51584 6016
rect 51520 5956 51524 6012
rect 51524 5956 51580 6012
rect 51580 5956 51584 6012
rect 51520 5952 51584 5956
rect 51600 6012 51664 6016
rect 51600 5956 51604 6012
rect 51604 5956 51660 6012
rect 51660 5956 51664 6012
rect 51600 5952 51664 5956
rect 51680 6012 51744 6016
rect 51680 5956 51684 6012
rect 51684 5956 51740 6012
rect 51740 5956 51744 6012
rect 51680 5952 51744 5956
rect 51760 6012 51824 6016
rect 51760 5956 51764 6012
rect 51764 5956 51820 6012
rect 51820 5956 51824 6012
rect 51760 5952 51824 5956
rect 15400 5468 15464 5472
rect 15400 5412 15404 5468
rect 15404 5412 15460 5468
rect 15460 5412 15464 5468
rect 15400 5408 15464 5412
rect 15480 5468 15544 5472
rect 15480 5412 15484 5468
rect 15484 5412 15540 5468
rect 15540 5412 15544 5468
rect 15480 5408 15544 5412
rect 15560 5468 15624 5472
rect 15560 5412 15564 5468
rect 15564 5412 15620 5468
rect 15620 5412 15624 5468
rect 15560 5408 15624 5412
rect 15640 5468 15704 5472
rect 15640 5412 15644 5468
rect 15644 5412 15700 5468
rect 15700 5412 15704 5468
rect 15640 5408 15704 5412
rect 29848 5468 29912 5472
rect 29848 5412 29852 5468
rect 29852 5412 29908 5468
rect 29908 5412 29912 5468
rect 29848 5408 29912 5412
rect 29928 5468 29992 5472
rect 29928 5412 29932 5468
rect 29932 5412 29988 5468
rect 29988 5412 29992 5468
rect 29928 5408 29992 5412
rect 30008 5468 30072 5472
rect 30008 5412 30012 5468
rect 30012 5412 30068 5468
rect 30068 5412 30072 5468
rect 30008 5408 30072 5412
rect 30088 5468 30152 5472
rect 30088 5412 30092 5468
rect 30092 5412 30148 5468
rect 30148 5412 30152 5468
rect 30088 5408 30152 5412
rect 44296 5468 44360 5472
rect 44296 5412 44300 5468
rect 44300 5412 44356 5468
rect 44356 5412 44360 5468
rect 44296 5408 44360 5412
rect 44376 5468 44440 5472
rect 44376 5412 44380 5468
rect 44380 5412 44436 5468
rect 44436 5412 44440 5468
rect 44376 5408 44440 5412
rect 44456 5468 44520 5472
rect 44456 5412 44460 5468
rect 44460 5412 44516 5468
rect 44516 5412 44520 5468
rect 44456 5408 44520 5412
rect 44536 5468 44600 5472
rect 44536 5412 44540 5468
rect 44540 5412 44596 5468
rect 44596 5412 44600 5468
rect 44536 5408 44600 5412
rect 8176 4924 8240 4928
rect 8176 4868 8180 4924
rect 8180 4868 8236 4924
rect 8236 4868 8240 4924
rect 8176 4864 8240 4868
rect 8256 4924 8320 4928
rect 8256 4868 8260 4924
rect 8260 4868 8316 4924
rect 8316 4868 8320 4924
rect 8256 4864 8320 4868
rect 8336 4924 8400 4928
rect 8336 4868 8340 4924
rect 8340 4868 8396 4924
rect 8396 4868 8400 4924
rect 8336 4864 8400 4868
rect 8416 4924 8480 4928
rect 8416 4868 8420 4924
rect 8420 4868 8476 4924
rect 8476 4868 8480 4924
rect 8416 4864 8480 4868
rect 22624 4924 22688 4928
rect 22624 4868 22628 4924
rect 22628 4868 22684 4924
rect 22684 4868 22688 4924
rect 22624 4864 22688 4868
rect 22704 4924 22768 4928
rect 22704 4868 22708 4924
rect 22708 4868 22764 4924
rect 22764 4868 22768 4924
rect 22704 4864 22768 4868
rect 22784 4924 22848 4928
rect 22784 4868 22788 4924
rect 22788 4868 22844 4924
rect 22844 4868 22848 4924
rect 22784 4864 22848 4868
rect 22864 4924 22928 4928
rect 22864 4868 22868 4924
rect 22868 4868 22924 4924
rect 22924 4868 22928 4924
rect 22864 4864 22928 4868
rect 37072 4924 37136 4928
rect 37072 4868 37076 4924
rect 37076 4868 37132 4924
rect 37132 4868 37136 4924
rect 37072 4864 37136 4868
rect 37152 4924 37216 4928
rect 37152 4868 37156 4924
rect 37156 4868 37212 4924
rect 37212 4868 37216 4924
rect 37152 4864 37216 4868
rect 37232 4924 37296 4928
rect 37232 4868 37236 4924
rect 37236 4868 37292 4924
rect 37292 4868 37296 4924
rect 37232 4864 37296 4868
rect 37312 4924 37376 4928
rect 37312 4868 37316 4924
rect 37316 4868 37372 4924
rect 37372 4868 37376 4924
rect 37312 4864 37376 4868
rect 51520 4924 51584 4928
rect 51520 4868 51524 4924
rect 51524 4868 51580 4924
rect 51580 4868 51584 4924
rect 51520 4864 51584 4868
rect 51600 4924 51664 4928
rect 51600 4868 51604 4924
rect 51604 4868 51660 4924
rect 51660 4868 51664 4924
rect 51600 4864 51664 4868
rect 51680 4924 51744 4928
rect 51680 4868 51684 4924
rect 51684 4868 51740 4924
rect 51740 4868 51744 4924
rect 51680 4864 51744 4868
rect 51760 4924 51824 4928
rect 51760 4868 51764 4924
rect 51764 4868 51820 4924
rect 51820 4868 51824 4924
rect 51760 4864 51824 4868
rect 15400 4380 15464 4384
rect 15400 4324 15404 4380
rect 15404 4324 15460 4380
rect 15460 4324 15464 4380
rect 15400 4320 15464 4324
rect 15480 4380 15544 4384
rect 15480 4324 15484 4380
rect 15484 4324 15540 4380
rect 15540 4324 15544 4380
rect 15480 4320 15544 4324
rect 15560 4380 15624 4384
rect 15560 4324 15564 4380
rect 15564 4324 15620 4380
rect 15620 4324 15624 4380
rect 15560 4320 15624 4324
rect 15640 4380 15704 4384
rect 15640 4324 15644 4380
rect 15644 4324 15700 4380
rect 15700 4324 15704 4380
rect 15640 4320 15704 4324
rect 29848 4380 29912 4384
rect 29848 4324 29852 4380
rect 29852 4324 29908 4380
rect 29908 4324 29912 4380
rect 29848 4320 29912 4324
rect 29928 4380 29992 4384
rect 29928 4324 29932 4380
rect 29932 4324 29988 4380
rect 29988 4324 29992 4380
rect 29928 4320 29992 4324
rect 30008 4380 30072 4384
rect 30008 4324 30012 4380
rect 30012 4324 30068 4380
rect 30068 4324 30072 4380
rect 30008 4320 30072 4324
rect 30088 4380 30152 4384
rect 30088 4324 30092 4380
rect 30092 4324 30148 4380
rect 30148 4324 30152 4380
rect 30088 4320 30152 4324
rect 44296 4380 44360 4384
rect 44296 4324 44300 4380
rect 44300 4324 44356 4380
rect 44356 4324 44360 4380
rect 44296 4320 44360 4324
rect 44376 4380 44440 4384
rect 44376 4324 44380 4380
rect 44380 4324 44436 4380
rect 44436 4324 44440 4380
rect 44376 4320 44440 4324
rect 44456 4380 44520 4384
rect 44456 4324 44460 4380
rect 44460 4324 44516 4380
rect 44516 4324 44520 4380
rect 44456 4320 44520 4324
rect 44536 4380 44600 4384
rect 44536 4324 44540 4380
rect 44540 4324 44596 4380
rect 44596 4324 44600 4380
rect 44536 4320 44600 4324
rect 8176 3836 8240 3840
rect 8176 3780 8180 3836
rect 8180 3780 8236 3836
rect 8236 3780 8240 3836
rect 8176 3776 8240 3780
rect 8256 3836 8320 3840
rect 8256 3780 8260 3836
rect 8260 3780 8316 3836
rect 8316 3780 8320 3836
rect 8256 3776 8320 3780
rect 8336 3836 8400 3840
rect 8336 3780 8340 3836
rect 8340 3780 8396 3836
rect 8396 3780 8400 3836
rect 8336 3776 8400 3780
rect 8416 3836 8480 3840
rect 8416 3780 8420 3836
rect 8420 3780 8476 3836
rect 8476 3780 8480 3836
rect 8416 3776 8480 3780
rect 22624 3836 22688 3840
rect 22624 3780 22628 3836
rect 22628 3780 22684 3836
rect 22684 3780 22688 3836
rect 22624 3776 22688 3780
rect 22704 3836 22768 3840
rect 22704 3780 22708 3836
rect 22708 3780 22764 3836
rect 22764 3780 22768 3836
rect 22704 3776 22768 3780
rect 22784 3836 22848 3840
rect 22784 3780 22788 3836
rect 22788 3780 22844 3836
rect 22844 3780 22848 3836
rect 22784 3776 22848 3780
rect 22864 3836 22928 3840
rect 22864 3780 22868 3836
rect 22868 3780 22924 3836
rect 22924 3780 22928 3836
rect 22864 3776 22928 3780
rect 37072 3836 37136 3840
rect 37072 3780 37076 3836
rect 37076 3780 37132 3836
rect 37132 3780 37136 3836
rect 37072 3776 37136 3780
rect 37152 3836 37216 3840
rect 37152 3780 37156 3836
rect 37156 3780 37212 3836
rect 37212 3780 37216 3836
rect 37152 3776 37216 3780
rect 37232 3836 37296 3840
rect 37232 3780 37236 3836
rect 37236 3780 37292 3836
rect 37292 3780 37296 3836
rect 37232 3776 37296 3780
rect 37312 3836 37376 3840
rect 37312 3780 37316 3836
rect 37316 3780 37372 3836
rect 37372 3780 37376 3836
rect 37312 3776 37376 3780
rect 51520 3836 51584 3840
rect 51520 3780 51524 3836
rect 51524 3780 51580 3836
rect 51580 3780 51584 3836
rect 51520 3776 51584 3780
rect 51600 3836 51664 3840
rect 51600 3780 51604 3836
rect 51604 3780 51660 3836
rect 51660 3780 51664 3836
rect 51600 3776 51664 3780
rect 51680 3836 51744 3840
rect 51680 3780 51684 3836
rect 51684 3780 51740 3836
rect 51740 3780 51744 3836
rect 51680 3776 51744 3780
rect 51760 3836 51824 3840
rect 51760 3780 51764 3836
rect 51764 3780 51820 3836
rect 51820 3780 51824 3836
rect 51760 3776 51824 3780
rect 15400 3292 15464 3296
rect 15400 3236 15404 3292
rect 15404 3236 15460 3292
rect 15460 3236 15464 3292
rect 15400 3232 15464 3236
rect 15480 3292 15544 3296
rect 15480 3236 15484 3292
rect 15484 3236 15540 3292
rect 15540 3236 15544 3292
rect 15480 3232 15544 3236
rect 15560 3292 15624 3296
rect 15560 3236 15564 3292
rect 15564 3236 15620 3292
rect 15620 3236 15624 3292
rect 15560 3232 15624 3236
rect 15640 3292 15704 3296
rect 15640 3236 15644 3292
rect 15644 3236 15700 3292
rect 15700 3236 15704 3292
rect 15640 3232 15704 3236
rect 29848 3292 29912 3296
rect 29848 3236 29852 3292
rect 29852 3236 29908 3292
rect 29908 3236 29912 3292
rect 29848 3232 29912 3236
rect 29928 3292 29992 3296
rect 29928 3236 29932 3292
rect 29932 3236 29988 3292
rect 29988 3236 29992 3292
rect 29928 3232 29992 3236
rect 30008 3292 30072 3296
rect 30008 3236 30012 3292
rect 30012 3236 30068 3292
rect 30068 3236 30072 3292
rect 30008 3232 30072 3236
rect 30088 3292 30152 3296
rect 30088 3236 30092 3292
rect 30092 3236 30148 3292
rect 30148 3236 30152 3292
rect 30088 3232 30152 3236
rect 44296 3292 44360 3296
rect 44296 3236 44300 3292
rect 44300 3236 44356 3292
rect 44356 3236 44360 3292
rect 44296 3232 44360 3236
rect 44376 3292 44440 3296
rect 44376 3236 44380 3292
rect 44380 3236 44436 3292
rect 44436 3236 44440 3292
rect 44376 3232 44440 3236
rect 44456 3292 44520 3296
rect 44456 3236 44460 3292
rect 44460 3236 44516 3292
rect 44516 3236 44520 3292
rect 44456 3232 44520 3236
rect 44536 3292 44600 3296
rect 44536 3236 44540 3292
rect 44540 3236 44596 3292
rect 44596 3236 44600 3292
rect 44536 3232 44600 3236
rect 8176 2748 8240 2752
rect 8176 2692 8180 2748
rect 8180 2692 8236 2748
rect 8236 2692 8240 2748
rect 8176 2688 8240 2692
rect 8256 2748 8320 2752
rect 8256 2692 8260 2748
rect 8260 2692 8316 2748
rect 8316 2692 8320 2748
rect 8256 2688 8320 2692
rect 8336 2748 8400 2752
rect 8336 2692 8340 2748
rect 8340 2692 8396 2748
rect 8396 2692 8400 2748
rect 8336 2688 8400 2692
rect 8416 2748 8480 2752
rect 8416 2692 8420 2748
rect 8420 2692 8476 2748
rect 8476 2692 8480 2748
rect 8416 2688 8480 2692
rect 22624 2748 22688 2752
rect 22624 2692 22628 2748
rect 22628 2692 22684 2748
rect 22684 2692 22688 2748
rect 22624 2688 22688 2692
rect 22704 2748 22768 2752
rect 22704 2692 22708 2748
rect 22708 2692 22764 2748
rect 22764 2692 22768 2748
rect 22704 2688 22768 2692
rect 22784 2748 22848 2752
rect 22784 2692 22788 2748
rect 22788 2692 22844 2748
rect 22844 2692 22848 2748
rect 22784 2688 22848 2692
rect 22864 2748 22928 2752
rect 22864 2692 22868 2748
rect 22868 2692 22924 2748
rect 22924 2692 22928 2748
rect 22864 2688 22928 2692
rect 37072 2748 37136 2752
rect 37072 2692 37076 2748
rect 37076 2692 37132 2748
rect 37132 2692 37136 2748
rect 37072 2688 37136 2692
rect 37152 2748 37216 2752
rect 37152 2692 37156 2748
rect 37156 2692 37212 2748
rect 37212 2692 37216 2748
rect 37152 2688 37216 2692
rect 37232 2748 37296 2752
rect 37232 2692 37236 2748
rect 37236 2692 37292 2748
rect 37292 2692 37296 2748
rect 37232 2688 37296 2692
rect 37312 2748 37376 2752
rect 37312 2692 37316 2748
rect 37316 2692 37372 2748
rect 37372 2692 37376 2748
rect 37312 2688 37376 2692
rect 51520 2748 51584 2752
rect 51520 2692 51524 2748
rect 51524 2692 51580 2748
rect 51580 2692 51584 2748
rect 51520 2688 51584 2692
rect 51600 2748 51664 2752
rect 51600 2692 51604 2748
rect 51604 2692 51660 2748
rect 51660 2692 51664 2748
rect 51600 2688 51664 2692
rect 51680 2748 51744 2752
rect 51680 2692 51684 2748
rect 51684 2692 51740 2748
rect 51740 2692 51744 2748
rect 51680 2688 51744 2692
rect 51760 2748 51824 2752
rect 51760 2692 51764 2748
rect 51764 2692 51820 2748
rect 51820 2692 51824 2748
rect 51760 2688 51824 2692
rect 15400 2204 15464 2208
rect 15400 2148 15404 2204
rect 15404 2148 15460 2204
rect 15460 2148 15464 2204
rect 15400 2144 15464 2148
rect 15480 2204 15544 2208
rect 15480 2148 15484 2204
rect 15484 2148 15540 2204
rect 15540 2148 15544 2204
rect 15480 2144 15544 2148
rect 15560 2204 15624 2208
rect 15560 2148 15564 2204
rect 15564 2148 15620 2204
rect 15620 2148 15624 2204
rect 15560 2144 15624 2148
rect 15640 2204 15704 2208
rect 15640 2148 15644 2204
rect 15644 2148 15700 2204
rect 15700 2148 15704 2204
rect 15640 2144 15704 2148
rect 29848 2204 29912 2208
rect 29848 2148 29852 2204
rect 29852 2148 29908 2204
rect 29908 2148 29912 2204
rect 29848 2144 29912 2148
rect 29928 2204 29992 2208
rect 29928 2148 29932 2204
rect 29932 2148 29988 2204
rect 29988 2148 29992 2204
rect 29928 2144 29992 2148
rect 30008 2204 30072 2208
rect 30008 2148 30012 2204
rect 30012 2148 30068 2204
rect 30068 2148 30072 2204
rect 30008 2144 30072 2148
rect 30088 2204 30152 2208
rect 30088 2148 30092 2204
rect 30092 2148 30148 2204
rect 30148 2148 30152 2204
rect 30088 2144 30152 2148
rect 44296 2204 44360 2208
rect 44296 2148 44300 2204
rect 44300 2148 44356 2204
rect 44356 2148 44360 2204
rect 44296 2144 44360 2148
rect 44376 2204 44440 2208
rect 44376 2148 44380 2204
rect 44380 2148 44436 2204
rect 44436 2148 44440 2204
rect 44376 2144 44440 2148
rect 44456 2204 44520 2208
rect 44456 2148 44460 2204
rect 44460 2148 44516 2204
rect 44516 2148 44520 2204
rect 44456 2144 44520 2148
rect 44536 2204 44600 2208
rect 44536 2148 44540 2204
rect 44540 2148 44596 2204
rect 44596 2148 44600 2204
rect 44536 2144 44600 2148
<< metal4 >>
rect 8168 33216 8488 33776
rect 8168 33152 8176 33216
rect 8240 33152 8256 33216
rect 8320 33152 8336 33216
rect 8400 33152 8416 33216
rect 8480 33152 8488 33216
rect 8168 32128 8488 33152
rect 8168 32064 8176 32128
rect 8240 32064 8256 32128
rect 8320 32064 8336 32128
rect 8400 32064 8416 32128
rect 8480 32064 8488 32128
rect 8168 31040 8488 32064
rect 8168 30976 8176 31040
rect 8240 30976 8256 31040
rect 8320 30976 8336 31040
rect 8400 30976 8416 31040
rect 8480 30976 8488 31040
rect 8168 29952 8488 30976
rect 8168 29888 8176 29952
rect 8240 29888 8256 29952
rect 8320 29888 8336 29952
rect 8400 29888 8416 29952
rect 8480 29888 8488 29952
rect 8168 28864 8488 29888
rect 8168 28800 8176 28864
rect 8240 28800 8256 28864
rect 8320 28800 8336 28864
rect 8400 28800 8416 28864
rect 8480 28800 8488 28864
rect 8168 27776 8488 28800
rect 8168 27712 8176 27776
rect 8240 27712 8256 27776
rect 8320 27712 8336 27776
rect 8400 27712 8416 27776
rect 8480 27712 8488 27776
rect 8168 26688 8488 27712
rect 8168 26624 8176 26688
rect 8240 26624 8256 26688
rect 8320 26624 8336 26688
rect 8400 26624 8416 26688
rect 8480 26624 8488 26688
rect 8168 25600 8488 26624
rect 8168 25536 8176 25600
rect 8240 25536 8256 25600
rect 8320 25536 8336 25600
rect 8400 25536 8416 25600
rect 8480 25536 8488 25600
rect 8168 24512 8488 25536
rect 8168 24448 8176 24512
rect 8240 24448 8256 24512
rect 8320 24448 8336 24512
rect 8400 24448 8416 24512
rect 8480 24448 8488 24512
rect 8168 23424 8488 24448
rect 8168 23360 8176 23424
rect 8240 23360 8256 23424
rect 8320 23360 8336 23424
rect 8400 23360 8416 23424
rect 8480 23360 8488 23424
rect 8168 22336 8488 23360
rect 8168 22272 8176 22336
rect 8240 22272 8256 22336
rect 8320 22272 8336 22336
rect 8400 22272 8416 22336
rect 8480 22272 8488 22336
rect 8168 21248 8488 22272
rect 8168 21184 8176 21248
rect 8240 21184 8256 21248
rect 8320 21184 8336 21248
rect 8400 21184 8416 21248
rect 8480 21184 8488 21248
rect 8168 20160 8488 21184
rect 8168 20096 8176 20160
rect 8240 20096 8256 20160
rect 8320 20096 8336 20160
rect 8400 20096 8416 20160
rect 8480 20096 8488 20160
rect 8168 19072 8488 20096
rect 8168 19008 8176 19072
rect 8240 19008 8256 19072
rect 8320 19008 8336 19072
rect 8400 19008 8416 19072
rect 8480 19008 8488 19072
rect 8168 17984 8488 19008
rect 8168 17920 8176 17984
rect 8240 17920 8256 17984
rect 8320 17920 8336 17984
rect 8400 17920 8416 17984
rect 8480 17920 8488 17984
rect 8168 16896 8488 17920
rect 8168 16832 8176 16896
rect 8240 16832 8256 16896
rect 8320 16832 8336 16896
rect 8400 16832 8416 16896
rect 8480 16832 8488 16896
rect 8168 15808 8488 16832
rect 8168 15744 8176 15808
rect 8240 15744 8256 15808
rect 8320 15744 8336 15808
rect 8400 15744 8416 15808
rect 8480 15744 8488 15808
rect 8168 14720 8488 15744
rect 8168 14656 8176 14720
rect 8240 14656 8256 14720
rect 8320 14656 8336 14720
rect 8400 14656 8416 14720
rect 8480 14656 8488 14720
rect 8168 13632 8488 14656
rect 8168 13568 8176 13632
rect 8240 13568 8256 13632
rect 8320 13568 8336 13632
rect 8400 13568 8416 13632
rect 8480 13568 8488 13632
rect 8168 12544 8488 13568
rect 8168 12480 8176 12544
rect 8240 12480 8256 12544
rect 8320 12480 8336 12544
rect 8400 12480 8416 12544
rect 8480 12480 8488 12544
rect 8168 11456 8488 12480
rect 8168 11392 8176 11456
rect 8240 11392 8256 11456
rect 8320 11392 8336 11456
rect 8400 11392 8416 11456
rect 8480 11392 8488 11456
rect 8168 10368 8488 11392
rect 8168 10304 8176 10368
rect 8240 10304 8256 10368
rect 8320 10304 8336 10368
rect 8400 10304 8416 10368
rect 8480 10304 8488 10368
rect 8168 9280 8488 10304
rect 8168 9216 8176 9280
rect 8240 9216 8256 9280
rect 8320 9216 8336 9280
rect 8400 9216 8416 9280
rect 8480 9216 8488 9280
rect 8168 8192 8488 9216
rect 8168 8128 8176 8192
rect 8240 8128 8256 8192
rect 8320 8128 8336 8192
rect 8400 8128 8416 8192
rect 8480 8128 8488 8192
rect 8168 7104 8488 8128
rect 8168 7040 8176 7104
rect 8240 7040 8256 7104
rect 8320 7040 8336 7104
rect 8400 7040 8416 7104
rect 8480 7040 8488 7104
rect 8168 6016 8488 7040
rect 8168 5952 8176 6016
rect 8240 5952 8256 6016
rect 8320 5952 8336 6016
rect 8400 5952 8416 6016
rect 8480 5952 8488 6016
rect 8168 4928 8488 5952
rect 8168 4864 8176 4928
rect 8240 4864 8256 4928
rect 8320 4864 8336 4928
rect 8400 4864 8416 4928
rect 8480 4864 8488 4928
rect 8168 3840 8488 4864
rect 8168 3776 8176 3840
rect 8240 3776 8256 3840
rect 8320 3776 8336 3840
rect 8400 3776 8416 3840
rect 8480 3776 8488 3840
rect 8168 2752 8488 3776
rect 8168 2688 8176 2752
rect 8240 2688 8256 2752
rect 8320 2688 8336 2752
rect 8400 2688 8416 2752
rect 8480 2688 8488 2752
rect 8168 2128 8488 2688
rect 15392 33760 15712 33776
rect 15392 33696 15400 33760
rect 15464 33696 15480 33760
rect 15544 33696 15560 33760
rect 15624 33696 15640 33760
rect 15704 33696 15712 33760
rect 15392 32672 15712 33696
rect 15392 32608 15400 32672
rect 15464 32608 15480 32672
rect 15544 32608 15560 32672
rect 15624 32608 15640 32672
rect 15704 32608 15712 32672
rect 15392 31584 15712 32608
rect 15392 31520 15400 31584
rect 15464 31520 15480 31584
rect 15544 31520 15560 31584
rect 15624 31520 15640 31584
rect 15704 31520 15712 31584
rect 15392 30496 15712 31520
rect 15392 30432 15400 30496
rect 15464 30432 15480 30496
rect 15544 30432 15560 30496
rect 15624 30432 15640 30496
rect 15704 30432 15712 30496
rect 15392 29408 15712 30432
rect 15392 29344 15400 29408
rect 15464 29344 15480 29408
rect 15544 29344 15560 29408
rect 15624 29344 15640 29408
rect 15704 29344 15712 29408
rect 15392 28320 15712 29344
rect 15392 28256 15400 28320
rect 15464 28256 15480 28320
rect 15544 28256 15560 28320
rect 15624 28256 15640 28320
rect 15704 28256 15712 28320
rect 15392 27232 15712 28256
rect 15392 27168 15400 27232
rect 15464 27168 15480 27232
rect 15544 27168 15560 27232
rect 15624 27168 15640 27232
rect 15704 27168 15712 27232
rect 15392 26144 15712 27168
rect 15392 26080 15400 26144
rect 15464 26080 15480 26144
rect 15544 26080 15560 26144
rect 15624 26080 15640 26144
rect 15704 26080 15712 26144
rect 15392 25056 15712 26080
rect 15392 24992 15400 25056
rect 15464 24992 15480 25056
rect 15544 24992 15560 25056
rect 15624 24992 15640 25056
rect 15704 24992 15712 25056
rect 15392 23968 15712 24992
rect 15392 23904 15400 23968
rect 15464 23904 15480 23968
rect 15544 23904 15560 23968
rect 15624 23904 15640 23968
rect 15704 23904 15712 23968
rect 15392 22880 15712 23904
rect 15392 22816 15400 22880
rect 15464 22816 15480 22880
rect 15544 22816 15560 22880
rect 15624 22816 15640 22880
rect 15704 22816 15712 22880
rect 15392 21792 15712 22816
rect 15392 21728 15400 21792
rect 15464 21728 15480 21792
rect 15544 21728 15560 21792
rect 15624 21728 15640 21792
rect 15704 21728 15712 21792
rect 15392 20704 15712 21728
rect 15392 20640 15400 20704
rect 15464 20640 15480 20704
rect 15544 20640 15560 20704
rect 15624 20640 15640 20704
rect 15704 20640 15712 20704
rect 15392 19616 15712 20640
rect 15392 19552 15400 19616
rect 15464 19552 15480 19616
rect 15544 19552 15560 19616
rect 15624 19552 15640 19616
rect 15704 19552 15712 19616
rect 15392 18528 15712 19552
rect 15392 18464 15400 18528
rect 15464 18464 15480 18528
rect 15544 18464 15560 18528
rect 15624 18464 15640 18528
rect 15704 18464 15712 18528
rect 15392 17440 15712 18464
rect 15392 17376 15400 17440
rect 15464 17376 15480 17440
rect 15544 17376 15560 17440
rect 15624 17376 15640 17440
rect 15704 17376 15712 17440
rect 15392 16352 15712 17376
rect 15392 16288 15400 16352
rect 15464 16288 15480 16352
rect 15544 16288 15560 16352
rect 15624 16288 15640 16352
rect 15704 16288 15712 16352
rect 15392 15264 15712 16288
rect 15392 15200 15400 15264
rect 15464 15200 15480 15264
rect 15544 15200 15560 15264
rect 15624 15200 15640 15264
rect 15704 15200 15712 15264
rect 15392 14176 15712 15200
rect 15392 14112 15400 14176
rect 15464 14112 15480 14176
rect 15544 14112 15560 14176
rect 15624 14112 15640 14176
rect 15704 14112 15712 14176
rect 15392 13088 15712 14112
rect 15392 13024 15400 13088
rect 15464 13024 15480 13088
rect 15544 13024 15560 13088
rect 15624 13024 15640 13088
rect 15704 13024 15712 13088
rect 15392 12000 15712 13024
rect 15392 11936 15400 12000
rect 15464 11936 15480 12000
rect 15544 11936 15560 12000
rect 15624 11936 15640 12000
rect 15704 11936 15712 12000
rect 15392 10912 15712 11936
rect 15392 10848 15400 10912
rect 15464 10848 15480 10912
rect 15544 10848 15560 10912
rect 15624 10848 15640 10912
rect 15704 10848 15712 10912
rect 15392 9824 15712 10848
rect 15392 9760 15400 9824
rect 15464 9760 15480 9824
rect 15544 9760 15560 9824
rect 15624 9760 15640 9824
rect 15704 9760 15712 9824
rect 15392 8736 15712 9760
rect 15392 8672 15400 8736
rect 15464 8672 15480 8736
rect 15544 8672 15560 8736
rect 15624 8672 15640 8736
rect 15704 8672 15712 8736
rect 15392 7648 15712 8672
rect 15392 7584 15400 7648
rect 15464 7584 15480 7648
rect 15544 7584 15560 7648
rect 15624 7584 15640 7648
rect 15704 7584 15712 7648
rect 15392 6560 15712 7584
rect 15392 6496 15400 6560
rect 15464 6496 15480 6560
rect 15544 6496 15560 6560
rect 15624 6496 15640 6560
rect 15704 6496 15712 6560
rect 15392 5472 15712 6496
rect 15392 5408 15400 5472
rect 15464 5408 15480 5472
rect 15544 5408 15560 5472
rect 15624 5408 15640 5472
rect 15704 5408 15712 5472
rect 15392 4384 15712 5408
rect 15392 4320 15400 4384
rect 15464 4320 15480 4384
rect 15544 4320 15560 4384
rect 15624 4320 15640 4384
rect 15704 4320 15712 4384
rect 15392 3296 15712 4320
rect 15392 3232 15400 3296
rect 15464 3232 15480 3296
rect 15544 3232 15560 3296
rect 15624 3232 15640 3296
rect 15704 3232 15712 3296
rect 15392 2208 15712 3232
rect 15392 2144 15400 2208
rect 15464 2144 15480 2208
rect 15544 2144 15560 2208
rect 15624 2144 15640 2208
rect 15704 2144 15712 2208
rect 15392 2128 15712 2144
rect 22616 33216 22936 33776
rect 22616 33152 22624 33216
rect 22688 33152 22704 33216
rect 22768 33152 22784 33216
rect 22848 33152 22864 33216
rect 22928 33152 22936 33216
rect 22616 32128 22936 33152
rect 22616 32064 22624 32128
rect 22688 32064 22704 32128
rect 22768 32064 22784 32128
rect 22848 32064 22864 32128
rect 22928 32064 22936 32128
rect 22616 31040 22936 32064
rect 22616 30976 22624 31040
rect 22688 30976 22704 31040
rect 22768 30976 22784 31040
rect 22848 30976 22864 31040
rect 22928 30976 22936 31040
rect 22616 29952 22936 30976
rect 22616 29888 22624 29952
rect 22688 29888 22704 29952
rect 22768 29888 22784 29952
rect 22848 29888 22864 29952
rect 22928 29888 22936 29952
rect 22616 28864 22936 29888
rect 22616 28800 22624 28864
rect 22688 28800 22704 28864
rect 22768 28800 22784 28864
rect 22848 28800 22864 28864
rect 22928 28800 22936 28864
rect 22616 27776 22936 28800
rect 22616 27712 22624 27776
rect 22688 27712 22704 27776
rect 22768 27712 22784 27776
rect 22848 27712 22864 27776
rect 22928 27712 22936 27776
rect 22616 26688 22936 27712
rect 22616 26624 22624 26688
rect 22688 26624 22704 26688
rect 22768 26624 22784 26688
rect 22848 26624 22864 26688
rect 22928 26624 22936 26688
rect 22616 25600 22936 26624
rect 22616 25536 22624 25600
rect 22688 25536 22704 25600
rect 22768 25536 22784 25600
rect 22848 25536 22864 25600
rect 22928 25536 22936 25600
rect 22616 24512 22936 25536
rect 22616 24448 22624 24512
rect 22688 24448 22704 24512
rect 22768 24448 22784 24512
rect 22848 24448 22864 24512
rect 22928 24448 22936 24512
rect 22616 23424 22936 24448
rect 22616 23360 22624 23424
rect 22688 23360 22704 23424
rect 22768 23360 22784 23424
rect 22848 23360 22864 23424
rect 22928 23360 22936 23424
rect 22616 22336 22936 23360
rect 22616 22272 22624 22336
rect 22688 22272 22704 22336
rect 22768 22272 22784 22336
rect 22848 22272 22864 22336
rect 22928 22272 22936 22336
rect 22616 21248 22936 22272
rect 22616 21184 22624 21248
rect 22688 21184 22704 21248
rect 22768 21184 22784 21248
rect 22848 21184 22864 21248
rect 22928 21184 22936 21248
rect 22616 20160 22936 21184
rect 22616 20096 22624 20160
rect 22688 20096 22704 20160
rect 22768 20096 22784 20160
rect 22848 20096 22864 20160
rect 22928 20096 22936 20160
rect 22616 19072 22936 20096
rect 22616 19008 22624 19072
rect 22688 19008 22704 19072
rect 22768 19008 22784 19072
rect 22848 19008 22864 19072
rect 22928 19008 22936 19072
rect 22616 17984 22936 19008
rect 22616 17920 22624 17984
rect 22688 17920 22704 17984
rect 22768 17920 22784 17984
rect 22848 17920 22864 17984
rect 22928 17920 22936 17984
rect 22616 16896 22936 17920
rect 22616 16832 22624 16896
rect 22688 16832 22704 16896
rect 22768 16832 22784 16896
rect 22848 16832 22864 16896
rect 22928 16832 22936 16896
rect 22616 15808 22936 16832
rect 22616 15744 22624 15808
rect 22688 15744 22704 15808
rect 22768 15744 22784 15808
rect 22848 15744 22864 15808
rect 22928 15744 22936 15808
rect 22616 14720 22936 15744
rect 22616 14656 22624 14720
rect 22688 14656 22704 14720
rect 22768 14656 22784 14720
rect 22848 14656 22864 14720
rect 22928 14656 22936 14720
rect 22616 13632 22936 14656
rect 22616 13568 22624 13632
rect 22688 13568 22704 13632
rect 22768 13568 22784 13632
rect 22848 13568 22864 13632
rect 22928 13568 22936 13632
rect 22616 12544 22936 13568
rect 22616 12480 22624 12544
rect 22688 12480 22704 12544
rect 22768 12480 22784 12544
rect 22848 12480 22864 12544
rect 22928 12480 22936 12544
rect 22616 11456 22936 12480
rect 22616 11392 22624 11456
rect 22688 11392 22704 11456
rect 22768 11392 22784 11456
rect 22848 11392 22864 11456
rect 22928 11392 22936 11456
rect 22616 10368 22936 11392
rect 22616 10304 22624 10368
rect 22688 10304 22704 10368
rect 22768 10304 22784 10368
rect 22848 10304 22864 10368
rect 22928 10304 22936 10368
rect 22616 9280 22936 10304
rect 22616 9216 22624 9280
rect 22688 9216 22704 9280
rect 22768 9216 22784 9280
rect 22848 9216 22864 9280
rect 22928 9216 22936 9280
rect 22616 8192 22936 9216
rect 22616 8128 22624 8192
rect 22688 8128 22704 8192
rect 22768 8128 22784 8192
rect 22848 8128 22864 8192
rect 22928 8128 22936 8192
rect 22616 7104 22936 8128
rect 22616 7040 22624 7104
rect 22688 7040 22704 7104
rect 22768 7040 22784 7104
rect 22848 7040 22864 7104
rect 22928 7040 22936 7104
rect 22616 6016 22936 7040
rect 22616 5952 22624 6016
rect 22688 5952 22704 6016
rect 22768 5952 22784 6016
rect 22848 5952 22864 6016
rect 22928 5952 22936 6016
rect 22616 4928 22936 5952
rect 22616 4864 22624 4928
rect 22688 4864 22704 4928
rect 22768 4864 22784 4928
rect 22848 4864 22864 4928
rect 22928 4864 22936 4928
rect 22616 3840 22936 4864
rect 22616 3776 22624 3840
rect 22688 3776 22704 3840
rect 22768 3776 22784 3840
rect 22848 3776 22864 3840
rect 22928 3776 22936 3840
rect 22616 2752 22936 3776
rect 22616 2688 22624 2752
rect 22688 2688 22704 2752
rect 22768 2688 22784 2752
rect 22848 2688 22864 2752
rect 22928 2688 22936 2752
rect 22616 2128 22936 2688
rect 29840 33760 30160 33776
rect 29840 33696 29848 33760
rect 29912 33696 29928 33760
rect 29992 33696 30008 33760
rect 30072 33696 30088 33760
rect 30152 33696 30160 33760
rect 29840 32672 30160 33696
rect 29840 32608 29848 32672
rect 29912 32608 29928 32672
rect 29992 32608 30008 32672
rect 30072 32608 30088 32672
rect 30152 32608 30160 32672
rect 29840 31584 30160 32608
rect 29840 31520 29848 31584
rect 29912 31520 29928 31584
rect 29992 31520 30008 31584
rect 30072 31520 30088 31584
rect 30152 31520 30160 31584
rect 29840 30496 30160 31520
rect 29840 30432 29848 30496
rect 29912 30432 29928 30496
rect 29992 30432 30008 30496
rect 30072 30432 30088 30496
rect 30152 30432 30160 30496
rect 29840 29408 30160 30432
rect 29840 29344 29848 29408
rect 29912 29344 29928 29408
rect 29992 29344 30008 29408
rect 30072 29344 30088 29408
rect 30152 29344 30160 29408
rect 29840 28320 30160 29344
rect 29840 28256 29848 28320
rect 29912 28256 29928 28320
rect 29992 28256 30008 28320
rect 30072 28256 30088 28320
rect 30152 28256 30160 28320
rect 29840 27232 30160 28256
rect 29840 27168 29848 27232
rect 29912 27168 29928 27232
rect 29992 27168 30008 27232
rect 30072 27168 30088 27232
rect 30152 27168 30160 27232
rect 29840 26144 30160 27168
rect 29840 26080 29848 26144
rect 29912 26080 29928 26144
rect 29992 26080 30008 26144
rect 30072 26080 30088 26144
rect 30152 26080 30160 26144
rect 29840 25056 30160 26080
rect 29840 24992 29848 25056
rect 29912 24992 29928 25056
rect 29992 24992 30008 25056
rect 30072 24992 30088 25056
rect 30152 24992 30160 25056
rect 29840 23968 30160 24992
rect 29840 23904 29848 23968
rect 29912 23904 29928 23968
rect 29992 23904 30008 23968
rect 30072 23904 30088 23968
rect 30152 23904 30160 23968
rect 29840 22880 30160 23904
rect 29840 22816 29848 22880
rect 29912 22816 29928 22880
rect 29992 22816 30008 22880
rect 30072 22816 30088 22880
rect 30152 22816 30160 22880
rect 29840 21792 30160 22816
rect 29840 21728 29848 21792
rect 29912 21728 29928 21792
rect 29992 21728 30008 21792
rect 30072 21728 30088 21792
rect 30152 21728 30160 21792
rect 29840 20704 30160 21728
rect 29840 20640 29848 20704
rect 29912 20640 29928 20704
rect 29992 20640 30008 20704
rect 30072 20640 30088 20704
rect 30152 20640 30160 20704
rect 29840 19616 30160 20640
rect 29840 19552 29848 19616
rect 29912 19552 29928 19616
rect 29992 19552 30008 19616
rect 30072 19552 30088 19616
rect 30152 19552 30160 19616
rect 29840 18528 30160 19552
rect 29840 18464 29848 18528
rect 29912 18464 29928 18528
rect 29992 18464 30008 18528
rect 30072 18464 30088 18528
rect 30152 18464 30160 18528
rect 29840 17440 30160 18464
rect 29840 17376 29848 17440
rect 29912 17376 29928 17440
rect 29992 17376 30008 17440
rect 30072 17376 30088 17440
rect 30152 17376 30160 17440
rect 29840 16352 30160 17376
rect 29840 16288 29848 16352
rect 29912 16288 29928 16352
rect 29992 16288 30008 16352
rect 30072 16288 30088 16352
rect 30152 16288 30160 16352
rect 29840 15264 30160 16288
rect 29840 15200 29848 15264
rect 29912 15200 29928 15264
rect 29992 15200 30008 15264
rect 30072 15200 30088 15264
rect 30152 15200 30160 15264
rect 29840 14176 30160 15200
rect 29840 14112 29848 14176
rect 29912 14112 29928 14176
rect 29992 14112 30008 14176
rect 30072 14112 30088 14176
rect 30152 14112 30160 14176
rect 29840 13088 30160 14112
rect 29840 13024 29848 13088
rect 29912 13024 29928 13088
rect 29992 13024 30008 13088
rect 30072 13024 30088 13088
rect 30152 13024 30160 13088
rect 29840 12000 30160 13024
rect 29840 11936 29848 12000
rect 29912 11936 29928 12000
rect 29992 11936 30008 12000
rect 30072 11936 30088 12000
rect 30152 11936 30160 12000
rect 29840 10912 30160 11936
rect 29840 10848 29848 10912
rect 29912 10848 29928 10912
rect 29992 10848 30008 10912
rect 30072 10848 30088 10912
rect 30152 10848 30160 10912
rect 29840 9824 30160 10848
rect 29840 9760 29848 9824
rect 29912 9760 29928 9824
rect 29992 9760 30008 9824
rect 30072 9760 30088 9824
rect 30152 9760 30160 9824
rect 29840 8736 30160 9760
rect 29840 8672 29848 8736
rect 29912 8672 29928 8736
rect 29992 8672 30008 8736
rect 30072 8672 30088 8736
rect 30152 8672 30160 8736
rect 29840 7648 30160 8672
rect 29840 7584 29848 7648
rect 29912 7584 29928 7648
rect 29992 7584 30008 7648
rect 30072 7584 30088 7648
rect 30152 7584 30160 7648
rect 29840 6560 30160 7584
rect 29840 6496 29848 6560
rect 29912 6496 29928 6560
rect 29992 6496 30008 6560
rect 30072 6496 30088 6560
rect 30152 6496 30160 6560
rect 29840 5472 30160 6496
rect 29840 5408 29848 5472
rect 29912 5408 29928 5472
rect 29992 5408 30008 5472
rect 30072 5408 30088 5472
rect 30152 5408 30160 5472
rect 29840 4384 30160 5408
rect 29840 4320 29848 4384
rect 29912 4320 29928 4384
rect 29992 4320 30008 4384
rect 30072 4320 30088 4384
rect 30152 4320 30160 4384
rect 29840 3296 30160 4320
rect 29840 3232 29848 3296
rect 29912 3232 29928 3296
rect 29992 3232 30008 3296
rect 30072 3232 30088 3296
rect 30152 3232 30160 3296
rect 29840 2208 30160 3232
rect 29840 2144 29848 2208
rect 29912 2144 29928 2208
rect 29992 2144 30008 2208
rect 30072 2144 30088 2208
rect 30152 2144 30160 2208
rect 29840 2128 30160 2144
rect 37064 33216 37384 33776
rect 37064 33152 37072 33216
rect 37136 33152 37152 33216
rect 37216 33152 37232 33216
rect 37296 33152 37312 33216
rect 37376 33152 37384 33216
rect 37064 32128 37384 33152
rect 37064 32064 37072 32128
rect 37136 32064 37152 32128
rect 37216 32064 37232 32128
rect 37296 32064 37312 32128
rect 37376 32064 37384 32128
rect 37064 31040 37384 32064
rect 37064 30976 37072 31040
rect 37136 30976 37152 31040
rect 37216 30976 37232 31040
rect 37296 30976 37312 31040
rect 37376 30976 37384 31040
rect 37064 29952 37384 30976
rect 37064 29888 37072 29952
rect 37136 29888 37152 29952
rect 37216 29888 37232 29952
rect 37296 29888 37312 29952
rect 37376 29888 37384 29952
rect 37064 28864 37384 29888
rect 37064 28800 37072 28864
rect 37136 28800 37152 28864
rect 37216 28800 37232 28864
rect 37296 28800 37312 28864
rect 37376 28800 37384 28864
rect 37064 27776 37384 28800
rect 37064 27712 37072 27776
rect 37136 27712 37152 27776
rect 37216 27712 37232 27776
rect 37296 27712 37312 27776
rect 37376 27712 37384 27776
rect 37064 26688 37384 27712
rect 37064 26624 37072 26688
rect 37136 26624 37152 26688
rect 37216 26624 37232 26688
rect 37296 26624 37312 26688
rect 37376 26624 37384 26688
rect 37064 25600 37384 26624
rect 37064 25536 37072 25600
rect 37136 25536 37152 25600
rect 37216 25536 37232 25600
rect 37296 25536 37312 25600
rect 37376 25536 37384 25600
rect 37064 24512 37384 25536
rect 37064 24448 37072 24512
rect 37136 24448 37152 24512
rect 37216 24448 37232 24512
rect 37296 24448 37312 24512
rect 37376 24448 37384 24512
rect 37064 23424 37384 24448
rect 37064 23360 37072 23424
rect 37136 23360 37152 23424
rect 37216 23360 37232 23424
rect 37296 23360 37312 23424
rect 37376 23360 37384 23424
rect 37064 22336 37384 23360
rect 37064 22272 37072 22336
rect 37136 22272 37152 22336
rect 37216 22272 37232 22336
rect 37296 22272 37312 22336
rect 37376 22272 37384 22336
rect 37064 21248 37384 22272
rect 37064 21184 37072 21248
rect 37136 21184 37152 21248
rect 37216 21184 37232 21248
rect 37296 21184 37312 21248
rect 37376 21184 37384 21248
rect 37064 20160 37384 21184
rect 37064 20096 37072 20160
rect 37136 20096 37152 20160
rect 37216 20096 37232 20160
rect 37296 20096 37312 20160
rect 37376 20096 37384 20160
rect 37064 19072 37384 20096
rect 37064 19008 37072 19072
rect 37136 19008 37152 19072
rect 37216 19008 37232 19072
rect 37296 19008 37312 19072
rect 37376 19008 37384 19072
rect 37064 17984 37384 19008
rect 37064 17920 37072 17984
rect 37136 17920 37152 17984
rect 37216 17920 37232 17984
rect 37296 17920 37312 17984
rect 37376 17920 37384 17984
rect 37064 16896 37384 17920
rect 37064 16832 37072 16896
rect 37136 16832 37152 16896
rect 37216 16832 37232 16896
rect 37296 16832 37312 16896
rect 37376 16832 37384 16896
rect 37064 15808 37384 16832
rect 37064 15744 37072 15808
rect 37136 15744 37152 15808
rect 37216 15744 37232 15808
rect 37296 15744 37312 15808
rect 37376 15744 37384 15808
rect 37064 14720 37384 15744
rect 37064 14656 37072 14720
rect 37136 14656 37152 14720
rect 37216 14656 37232 14720
rect 37296 14656 37312 14720
rect 37376 14656 37384 14720
rect 37064 13632 37384 14656
rect 37064 13568 37072 13632
rect 37136 13568 37152 13632
rect 37216 13568 37232 13632
rect 37296 13568 37312 13632
rect 37376 13568 37384 13632
rect 37064 12544 37384 13568
rect 37064 12480 37072 12544
rect 37136 12480 37152 12544
rect 37216 12480 37232 12544
rect 37296 12480 37312 12544
rect 37376 12480 37384 12544
rect 37064 11456 37384 12480
rect 37064 11392 37072 11456
rect 37136 11392 37152 11456
rect 37216 11392 37232 11456
rect 37296 11392 37312 11456
rect 37376 11392 37384 11456
rect 37064 10368 37384 11392
rect 37064 10304 37072 10368
rect 37136 10304 37152 10368
rect 37216 10304 37232 10368
rect 37296 10304 37312 10368
rect 37376 10304 37384 10368
rect 37064 9280 37384 10304
rect 37064 9216 37072 9280
rect 37136 9216 37152 9280
rect 37216 9216 37232 9280
rect 37296 9216 37312 9280
rect 37376 9216 37384 9280
rect 37064 8192 37384 9216
rect 37064 8128 37072 8192
rect 37136 8128 37152 8192
rect 37216 8128 37232 8192
rect 37296 8128 37312 8192
rect 37376 8128 37384 8192
rect 37064 7104 37384 8128
rect 37064 7040 37072 7104
rect 37136 7040 37152 7104
rect 37216 7040 37232 7104
rect 37296 7040 37312 7104
rect 37376 7040 37384 7104
rect 37064 6016 37384 7040
rect 37064 5952 37072 6016
rect 37136 5952 37152 6016
rect 37216 5952 37232 6016
rect 37296 5952 37312 6016
rect 37376 5952 37384 6016
rect 37064 4928 37384 5952
rect 37064 4864 37072 4928
rect 37136 4864 37152 4928
rect 37216 4864 37232 4928
rect 37296 4864 37312 4928
rect 37376 4864 37384 4928
rect 37064 3840 37384 4864
rect 37064 3776 37072 3840
rect 37136 3776 37152 3840
rect 37216 3776 37232 3840
rect 37296 3776 37312 3840
rect 37376 3776 37384 3840
rect 37064 2752 37384 3776
rect 37064 2688 37072 2752
rect 37136 2688 37152 2752
rect 37216 2688 37232 2752
rect 37296 2688 37312 2752
rect 37376 2688 37384 2752
rect 37064 2128 37384 2688
rect 44288 33760 44608 33776
rect 44288 33696 44296 33760
rect 44360 33696 44376 33760
rect 44440 33696 44456 33760
rect 44520 33696 44536 33760
rect 44600 33696 44608 33760
rect 44288 32672 44608 33696
rect 44288 32608 44296 32672
rect 44360 32608 44376 32672
rect 44440 32608 44456 32672
rect 44520 32608 44536 32672
rect 44600 32608 44608 32672
rect 44288 31584 44608 32608
rect 44288 31520 44296 31584
rect 44360 31520 44376 31584
rect 44440 31520 44456 31584
rect 44520 31520 44536 31584
rect 44600 31520 44608 31584
rect 44288 30496 44608 31520
rect 44288 30432 44296 30496
rect 44360 30432 44376 30496
rect 44440 30432 44456 30496
rect 44520 30432 44536 30496
rect 44600 30432 44608 30496
rect 44288 29408 44608 30432
rect 44288 29344 44296 29408
rect 44360 29344 44376 29408
rect 44440 29344 44456 29408
rect 44520 29344 44536 29408
rect 44600 29344 44608 29408
rect 44288 28320 44608 29344
rect 44288 28256 44296 28320
rect 44360 28256 44376 28320
rect 44440 28256 44456 28320
rect 44520 28256 44536 28320
rect 44600 28256 44608 28320
rect 44288 27232 44608 28256
rect 44288 27168 44296 27232
rect 44360 27168 44376 27232
rect 44440 27168 44456 27232
rect 44520 27168 44536 27232
rect 44600 27168 44608 27232
rect 44288 26144 44608 27168
rect 44288 26080 44296 26144
rect 44360 26080 44376 26144
rect 44440 26080 44456 26144
rect 44520 26080 44536 26144
rect 44600 26080 44608 26144
rect 44288 25056 44608 26080
rect 44288 24992 44296 25056
rect 44360 24992 44376 25056
rect 44440 24992 44456 25056
rect 44520 24992 44536 25056
rect 44600 24992 44608 25056
rect 44288 23968 44608 24992
rect 44288 23904 44296 23968
rect 44360 23904 44376 23968
rect 44440 23904 44456 23968
rect 44520 23904 44536 23968
rect 44600 23904 44608 23968
rect 44288 22880 44608 23904
rect 44288 22816 44296 22880
rect 44360 22816 44376 22880
rect 44440 22816 44456 22880
rect 44520 22816 44536 22880
rect 44600 22816 44608 22880
rect 44288 21792 44608 22816
rect 44288 21728 44296 21792
rect 44360 21728 44376 21792
rect 44440 21728 44456 21792
rect 44520 21728 44536 21792
rect 44600 21728 44608 21792
rect 44288 20704 44608 21728
rect 44288 20640 44296 20704
rect 44360 20640 44376 20704
rect 44440 20640 44456 20704
rect 44520 20640 44536 20704
rect 44600 20640 44608 20704
rect 44288 19616 44608 20640
rect 44288 19552 44296 19616
rect 44360 19552 44376 19616
rect 44440 19552 44456 19616
rect 44520 19552 44536 19616
rect 44600 19552 44608 19616
rect 44288 18528 44608 19552
rect 44288 18464 44296 18528
rect 44360 18464 44376 18528
rect 44440 18464 44456 18528
rect 44520 18464 44536 18528
rect 44600 18464 44608 18528
rect 44288 17440 44608 18464
rect 44288 17376 44296 17440
rect 44360 17376 44376 17440
rect 44440 17376 44456 17440
rect 44520 17376 44536 17440
rect 44600 17376 44608 17440
rect 44288 16352 44608 17376
rect 44288 16288 44296 16352
rect 44360 16288 44376 16352
rect 44440 16288 44456 16352
rect 44520 16288 44536 16352
rect 44600 16288 44608 16352
rect 44288 15264 44608 16288
rect 44288 15200 44296 15264
rect 44360 15200 44376 15264
rect 44440 15200 44456 15264
rect 44520 15200 44536 15264
rect 44600 15200 44608 15264
rect 44288 14176 44608 15200
rect 44288 14112 44296 14176
rect 44360 14112 44376 14176
rect 44440 14112 44456 14176
rect 44520 14112 44536 14176
rect 44600 14112 44608 14176
rect 44288 13088 44608 14112
rect 44288 13024 44296 13088
rect 44360 13024 44376 13088
rect 44440 13024 44456 13088
rect 44520 13024 44536 13088
rect 44600 13024 44608 13088
rect 44288 12000 44608 13024
rect 44288 11936 44296 12000
rect 44360 11936 44376 12000
rect 44440 11936 44456 12000
rect 44520 11936 44536 12000
rect 44600 11936 44608 12000
rect 44288 10912 44608 11936
rect 44288 10848 44296 10912
rect 44360 10848 44376 10912
rect 44440 10848 44456 10912
rect 44520 10848 44536 10912
rect 44600 10848 44608 10912
rect 44288 9824 44608 10848
rect 44288 9760 44296 9824
rect 44360 9760 44376 9824
rect 44440 9760 44456 9824
rect 44520 9760 44536 9824
rect 44600 9760 44608 9824
rect 44288 8736 44608 9760
rect 44288 8672 44296 8736
rect 44360 8672 44376 8736
rect 44440 8672 44456 8736
rect 44520 8672 44536 8736
rect 44600 8672 44608 8736
rect 44288 7648 44608 8672
rect 44288 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44536 7648
rect 44600 7584 44608 7648
rect 44288 6560 44608 7584
rect 44288 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44536 6560
rect 44600 6496 44608 6560
rect 44288 5472 44608 6496
rect 44288 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44536 5472
rect 44600 5408 44608 5472
rect 44288 4384 44608 5408
rect 44288 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44536 4384
rect 44600 4320 44608 4384
rect 44288 3296 44608 4320
rect 44288 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44536 3296
rect 44600 3232 44608 3296
rect 44288 2208 44608 3232
rect 44288 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44536 2208
rect 44600 2144 44608 2208
rect 44288 2128 44608 2144
rect 51512 33216 51832 33776
rect 51512 33152 51520 33216
rect 51584 33152 51600 33216
rect 51664 33152 51680 33216
rect 51744 33152 51760 33216
rect 51824 33152 51832 33216
rect 51512 32128 51832 33152
rect 51512 32064 51520 32128
rect 51584 32064 51600 32128
rect 51664 32064 51680 32128
rect 51744 32064 51760 32128
rect 51824 32064 51832 32128
rect 51512 31040 51832 32064
rect 51512 30976 51520 31040
rect 51584 30976 51600 31040
rect 51664 30976 51680 31040
rect 51744 30976 51760 31040
rect 51824 30976 51832 31040
rect 51512 29952 51832 30976
rect 51512 29888 51520 29952
rect 51584 29888 51600 29952
rect 51664 29888 51680 29952
rect 51744 29888 51760 29952
rect 51824 29888 51832 29952
rect 51512 28864 51832 29888
rect 51512 28800 51520 28864
rect 51584 28800 51600 28864
rect 51664 28800 51680 28864
rect 51744 28800 51760 28864
rect 51824 28800 51832 28864
rect 51512 27776 51832 28800
rect 51512 27712 51520 27776
rect 51584 27712 51600 27776
rect 51664 27712 51680 27776
rect 51744 27712 51760 27776
rect 51824 27712 51832 27776
rect 51512 26688 51832 27712
rect 51512 26624 51520 26688
rect 51584 26624 51600 26688
rect 51664 26624 51680 26688
rect 51744 26624 51760 26688
rect 51824 26624 51832 26688
rect 51512 25600 51832 26624
rect 51512 25536 51520 25600
rect 51584 25536 51600 25600
rect 51664 25536 51680 25600
rect 51744 25536 51760 25600
rect 51824 25536 51832 25600
rect 51512 24512 51832 25536
rect 51512 24448 51520 24512
rect 51584 24448 51600 24512
rect 51664 24448 51680 24512
rect 51744 24448 51760 24512
rect 51824 24448 51832 24512
rect 51512 23424 51832 24448
rect 51512 23360 51520 23424
rect 51584 23360 51600 23424
rect 51664 23360 51680 23424
rect 51744 23360 51760 23424
rect 51824 23360 51832 23424
rect 51512 22336 51832 23360
rect 51512 22272 51520 22336
rect 51584 22272 51600 22336
rect 51664 22272 51680 22336
rect 51744 22272 51760 22336
rect 51824 22272 51832 22336
rect 51512 21248 51832 22272
rect 51512 21184 51520 21248
rect 51584 21184 51600 21248
rect 51664 21184 51680 21248
rect 51744 21184 51760 21248
rect 51824 21184 51832 21248
rect 51512 20160 51832 21184
rect 51512 20096 51520 20160
rect 51584 20096 51600 20160
rect 51664 20096 51680 20160
rect 51744 20096 51760 20160
rect 51824 20096 51832 20160
rect 51512 19072 51832 20096
rect 51512 19008 51520 19072
rect 51584 19008 51600 19072
rect 51664 19008 51680 19072
rect 51744 19008 51760 19072
rect 51824 19008 51832 19072
rect 51512 17984 51832 19008
rect 51512 17920 51520 17984
rect 51584 17920 51600 17984
rect 51664 17920 51680 17984
rect 51744 17920 51760 17984
rect 51824 17920 51832 17984
rect 51512 16896 51832 17920
rect 51512 16832 51520 16896
rect 51584 16832 51600 16896
rect 51664 16832 51680 16896
rect 51744 16832 51760 16896
rect 51824 16832 51832 16896
rect 51512 15808 51832 16832
rect 51512 15744 51520 15808
rect 51584 15744 51600 15808
rect 51664 15744 51680 15808
rect 51744 15744 51760 15808
rect 51824 15744 51832 15808
rect 51512 14720 51832 15744
rect 51512 14656 51520 14720
rect 51584 14656 51600 14720
rect 51664 14656 51680 14720
rect 51744 14656 51760 14720
rect 51824 14656 51832 14720
rect 51512 13632 51832 14656
rect 51512 13568 51520 13632
rect 51584 13568 51600 13632
rect 51664 13568 51680 13632
rect 51744 13568 51760 13632
rect 51824 13568 51832 13632
rect 51512 12544 51832 13568
rect 51512 12480 51520 12544
rect 51584 12480 51600 12544
rect 51664 12480 51680 12544
rect 51744 12480 51760 12544
rect 51824 12480 51832 12544
rect 51512 11456 51832 12480
rect 51512 11392 51520 11456
rect 51584 11392 51600 11456
rect 51664 11392 51680 11456
rect 51744 11392 51760 11456
rect 51824 11392 51832 11456
rect 51512 10368 51832 11392
rect 51512 10304 51520 10368
rect 51584 10304 51600 10368
rect 51664 10304 51680 10368
rect 51744 10304 51760 10368
rect 51824 10304 51832 10368
rect 51512 9280 51832 10304
rect 51512 9216 51520 9280
rect 51584 9216 51600 9280
rect 51664 9216 51680 9280
rect 51744 9216 51760 9280
rect 51824 9216 51832 9280
rect 51512 8192 51832 9216
rect 51512 8128 51520 8192
rect 51584 8128 51600 8192
rect 51664 8128 51680 8192
rect 51744 8128 51760 8192
rect 51824 8128 51832 8192
rect 51512 7104 51832 8128
rect 51512 7040 51520 7104
rect 51584 7040 51600 7104
rect 51664 7040 51680 7104
rect 51744 7040 51760 7104
rect 51824 7040 51832 7104
rect 51512 6016 51832 7040
rect 51512 5952 51520 6016
rect 51584 5952 51600 6016
rect 51664 5952 51680 6016
rect 51744 5952 51760 6016
rect 51824 5952 51832 6016
rect 51512 4928 51832 5952
rect 51512 4864 51520 4928
rect 51584 4864 51600 4928
rect 51664 4864 51680 4928
rect 51744 4864 51760 4928
rect 51824 4864 51832 4928
rect 51512 3840 51832 4864
rect 51512 3776 51520 3840
rect 51584 3776 51600 3840
rect 51664 3776 51680 3840
rect 51744 3776 51760 3840
rect 51824 3776 51832 3840
rect 51512 2752 51832 3776
rect 51512 2688 51520 2752
rect 51584 2688 51600 2752
rect 51664 2688 51680 2752
rect 51744 2688 51760 2752
rect 51824 2688 51832 2752
rect 51512 2128 51832 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__0485__1_A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 33764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1649977179
transform -1 0 21712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__A
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__A
timestamp 1649977179
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1649977179
transform -1 0 14628 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__B
timestamp 1649977179
transform -1 0 15640 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A
timestamp 1649977179
transform 1 0 18124 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1649977179
transform 1 0 2944 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A
timestamp 1649977179
transform -1 0 2576 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A
timestamp 1649977179
transform -1 0 4600 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__C
timestamp 1649977179
transform -1 0 6256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 1649977179
transform -1 0 20056 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A1
timestamp 1649977179
transform -1 0 23092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__C
timestamp 1649977179
transform 1 0 24932 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__A
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__B
timestamp 1649977179
transform -1 0 24564 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A
timestamp 1649977179
transform 1 0 16744 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1649977179
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A
timestamp 1649977179
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__B
timestamp 1649977179
transform -1 0 21344 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A
timestamp 1649977179
transform 1 0 27324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1649977179
transform 1 0 26312 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__A
timestamp 1649977179
transform -1 0 23368 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__B
timestamp 1649977179
transform -1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__C
timestamp 1649977179
transform -1 0 21344 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 1649977179
transform 1 0 19596 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B
timestamp 1649977179
transform -1 0 40296 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__D
timestamp 1649977179
transform 1 0 27508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1649977179
transform -1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A
timestamp 1649977179
transform -1 0 56120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A
timestamp 1649977179
transform 1 0 53728 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1649977179
transform -1 0 45172 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1649977179
transform 1 0 46276 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 1649977179
transform -1 0 43700 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A
timestamp 1649977179
transform 1 0 50876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A
timestamp 1649977179
transform 1 0 44160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1649977179
transform 1 0 45264 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1649977179
transform -1 0 50324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__C1
timestamp 1649977179
transform -1 0 49864 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B
timestamp 1649977179
transform -1 0 54832 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__B1
timestamp 1649977179
transform 1 0 52072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B1
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B1
timestamp 1649977179
transform 1 0 47656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__C1
timestamp 1649977179
transform -1 0 47380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1649977179
transform 1 0 48208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B
timestamp 1649977179
transform -1 0 21344 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A_N
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1649977179
transform -1 0 32844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__B
timestamp 1649977179
transform 1 0 33212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__B
timestamp 1649977179
transform -1 0 41216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__C
timestamp 1649977179
transform 1 0 31464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__B1
timestamp 1649977179
transform -1 0 39744 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B1
timestamp 1649977179
transform 1 0 33120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__B1
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B1
timestamp 1649977179
transform 1 0 33304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A
timestamp 1649977179
transform -1 0 28152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B1
timestamp 1649977179
transform 1 0 33396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1649977179
transform -1 0 28060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A_N
timestamp 1649977179
transform 1 0 28888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__B1
timestamp 1649977179
transform 1 0 32108 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A2
timestamp 1649977179
transform -1 0 27508 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1649977179
transform -1 0 25852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1649977179
transform -1 0 27048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B1
timestamp 1649977179
transform -1 0 34132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1649977179
transform -1 0 36800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1649977179
transform 1 0 43424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__C1
timestamp 1649977179
transform 1 0 39192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B
timestamp 1649977179
transform -1 0 44436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A
timestamp 1649977179
transform -1 0 29992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B1
timestamp 1649977179
transform -1 0 34868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1649977179
transform 1 0 36616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B1
timestamp 1649977179
transform 1 0 35696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1649977179
transform -1 0 47196 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1649977179
transform -1 0 45724 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__B1
timestamp 1649977179
transform 1 0 46184 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1649977179
transform -1 0 46276 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B1
timestamp 1649977179
transform -1 0 46644 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1649977179
transform 1 0 32200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__C1
timestamp 1649977179
transform -1 0 29900 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A
timestamp 1649977179
transform -1 0 39376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__B
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A
timestamp 1649977179
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__B1
timestamp 1649977179
transform 1 0 22080 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__C1
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1649977179
transform -1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1649977179
transform 1 0 37444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A
timestamp 1649977179
transform 1 0 26864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1649977179
transform 1 0 32752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1649977179
transform 1 0 40112 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A
timestamp 1649977179
transform -1 0 42872 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__B
timestamp 1649977179
transform -1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__B
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A
timestamp 1649977179
transform 1 0 21160 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__B
timestamp 1649977179
transform 1 0 23736 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__B
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A
timestamp 1649977179
transform 1 0 15088 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__B
timestamp 1649977179
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__B
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B
timestamp 1649977179
transform -1 0 3128 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A
timestamp 1649977179
transform 1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__B
timestamp 1649977179
transform -1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1649977179
transform -1 0 1656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__B
timestamp 1649977179
transform -1 0 1656 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B
timestamp 1649977179
transform -1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A
timestamp 1649977179
transform -1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A
timestamp 1649977179
transform -1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B
timestamp 1649977179
transform -1 0 5336 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A
timestamp 1649977179
transform -1 0 15180 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__B
timestamp 1649977179
transform -1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__CLK
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__CLK
timestamp 1649977179
transform 1 0 3128 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__CLK
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__CLK
timestamp 1649977179
transform 1 0 3128 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__CLK
timestamp 1649977179
transform 1 0 9200 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__CLK
timestamp 1649977179
transform 1 0 17296 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__CLK
timestamp 1649977179
transform 1 0 24104 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__CLK
timestamp 1649977179
transform 1 0 18584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__CLK
timestamp 1649977179
transform 1 0 29348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__CLK
timestamp 1649977179
transform 1 0 23736 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__CLK
timestamp 1649977179
transform -1 0 3680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__CLK
timestamp 1649977179
transform -1 0 19596 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__CLK
timestamp 1649977179
transform 1 0 31188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__CLK
timestamp 1649977179
transform 1 0 32016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__CLK
timestamp 1649977179
transform -1 0 30820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__CLK
timestamp 1649977179
transform 1 0 30360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__CLK
timestamp 1649977179
transform -1 0 39376 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__CLK
timestamp 1649977179
transform -1 0 41952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__CLK
timestamp 1649977179
transform -1 0 7544 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__D
timestamp 1649977179
transform 1 0 9476 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__CLK
timestamp 1649977179
transform -1 0 1932 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__D
timestamp 1649977179
transform 1 0 4140 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__CLK
timestamp 1649977179
transform 1 0 1932 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__CLK
timestamp 1649977179
transform 1 0 3128 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__CLK
timestamp 1649977179
transform -1 0 55936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__D
timestamp 1649977179
transform -1 0 58236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__CLK
timestamp 1649977179
transform 1 0 55292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__CLK
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__D
timestamp 1649977179
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__CLK
timestamp 1649977179
transform 1 0 17848 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__CLK
timestamp 1649977179
transform -1 0 39376 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__CLK
timestamp 1649977179
transform 1 0 33856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__RESET_B
timestamp 1649977179
transform 1 0 5152 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__RESET_B
timestamp 1649977179
transform 1 0 3220 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__RESET_B
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__CLK
timestamp 1649977179
transform 1 0 18032 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__RESET_B
timestamp 1649977179
transform 1 0 18584 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__RESET_B
timestamp 1649977179
transform -1 0 29716 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__CLK
timestamp 1649977179
transform 1 0 24104 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__RESET_B
timestamp 1649977179
transform -1 0 26496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__RESET_B
timestamp 1649977179
transform 1 0 15640 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__CLK
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__RESET_B
timestamp 1649977179
transform 1 0 18584 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__CLK
timestamp 1649977179
transform 1 0 17572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__CLK
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__CLK
timestamp 1649977179
transform 1 0 26036 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__CLK
timestamp 1649977179
transform -1 0 5888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__CLK
timestamp 1649977179
transform -1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__CLK
timestamp 1649977179
transform -1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__CLK
timestamp 1649977179
transform -1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__CLK
timestamp 1649977179
transform 1 0 16100 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__CLK
timestamp 1649977179
transform -1 0 17020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__CLK
timestamp 1649977179
transform -1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__CLK
timestamp 1649977179
transform -1 0 26404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__CLK
timestamp 1649977179
transform 1 0 14720 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__CLK
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__CLK
timestamp 1649977179
transform 1 0 15456 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__CLK
timestamp 1649977179
transform -1 0 25852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__CLK
timestamp 1649977179
transform -1 0 32936 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__CLK
timestamp 1649977179
transform -1 0 37444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__D
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__CLK
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__D
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__CLK
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__CLK
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__CLK
timestamp 1649977179
transform 1 0 29072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__D
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__CLK
timestamp 1649977179
transform 1 0 25300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__CLK
timestamp 1649977179
transform 1 0 27600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A
timestamp 1649977179
transform -1 0 37720 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__A
timestamp 1649977179
transform 1 0 18584 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__A
timestamp 1649977179
transform 1 0 4600 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__A
timestamp 1649977179
transform -1 0 57408 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__A
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__A
timestamp 1649977179
transform 1 0 57224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__A
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A
timestamp 1649977179
transform 1 0 25024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__A
timestamp 1649977179
transform -1 0 16928 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__A
timestamp 1649977179
transform -1 0 50416 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__A
timestamp 1649977179
transform -1 0 49496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__A
timestamp 1649977179
transform -1 0 46644 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__A
timestamp 1649977179
transform -1 0 33120 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A
timestamp 1649977179
transform -1 0 28704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A
timestamp 1649977179
transform -1 0 2024 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A
timestamp 1649977179
transform -1 0 23552 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_master_A
timestamp 1649977179
transform -1 0 18308 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_clk_master_A
timestamp 1649977179
transform 1 0 12512 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_clk_master_A
timestamp 1649977179
transform -1 0 12420 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_clk_master_A
timestamp 1649977179
transform 1 0 27416 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_clk_master_A
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 44068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 57592 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 58236 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 25208 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 53084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 1748 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 28060 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 57500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_net99_2_A
timestamp 1649977179
transform -1 0 34040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_A
timestamp 1649977179
transform 1 0 25116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output26_A
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_A
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output29_A
timestamp 1649977179
transform -1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 1649977179
transform 1 0 52716 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater79_A
timestamp 1649977179
transform 1 0 18676 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater84_A
timestamp 1649977179
transform -1 0 16192 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater93_A
timestamp 1649977179
transform -1 0 43884 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater94_A
timestamp 1649977179
transform -1 0 44804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 6992 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 4600 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 6808 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 4600 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 5704 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 4048 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 8004 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 8096 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 9476 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1649977179
transform -1 0 6808 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N
timestamp 1649977179
transform -1 0 7360 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 7544 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 4048 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 9476 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 3404 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 3036 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 35512 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 34960 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 35696 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 36248 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 34960 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 35328 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
timestamp 1649977179
transform -1 0 34224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1649977179
transform -1 0 39100 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_GATE_N
timestamp 1649977179
transform -1 0 39652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf_TE_B
timestamp 1649977179
transform 1 0 31188 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 37352 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 37904 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 38548 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 39100 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 35512 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 35880 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf_TE_B
timestamp 1649977179
transform -1 0 29072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1649977179
transform -1 0 35696 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_GATE_N
timestamp 1649977179
transform -1 0 36064 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 34684 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 34040 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf_A
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 34592 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_GATE_N
timestamp 1649977179
transform 1 0 34960 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf_A
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.ro_block_I.ro_pol.tribuf.t_buf_TE_B
timestamp 1649977179
transform -1 0 27968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_w0.ro_block_I.ro_pol_eve.tribuf.t_buf_TE_B
timestamp 1649977179
transform -1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 46000 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 46552 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 46644 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
timestamp 1649977179
transform -1 0 47748 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 51336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 46644 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 50784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn_D
timestamp 1649977179
transform -1 0 47748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn_D
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf_TE_B
timestamp 1649977179
transform -1 0 48760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.ro_block_I.ro_pol.tribuf.t_buf_TE_B
timestamp 1649977179
transform -1 0 21804 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wrapper_cell_loop\[0\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf_TE_B
timestamp 1649977179
transform -1 0 19688 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42
timestamp 1649977179
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1649977179
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_147
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_203
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1649977179
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_263
timestamp 1649977179
transform 1 0 25300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1649977179
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1649977179
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1649977179
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_313
timestamp 1649977179
transform 1 0 29900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_325
timestamp 1649977179
transform 1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1649977179
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1649977179
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1649977179
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_401
timestamp 1649977179
transform 1 0 37996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_405
timestamp 1649977179
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_413 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39100 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1649977179
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1649977179
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1649977179
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_449
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_457
timestamp 1649977179
transform 1 0 43148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1649977179
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_467
timestamp 1649977179
transform 1 0 44068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1649977179
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1649977179
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1649977179
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_505
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_513
timestamp 1649977179
transform 1 0 48300 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_518
timestamp 1649977179
transform 1 0 48760 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1649977179
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_545
timestamp 1649977179
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1649977179
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_561
timestamp 1649977179
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_569
timestamp 1649977179
transform 1 0 53452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_581
timestamp 1649977179
transform 1 0 54556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1649977179
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1649977179
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_601
timestamp 1649977179
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_613
timestamp 1649977179
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1649977179
transform 1 0 58236 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_143
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_155
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_216
timestamp 1649977179
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_289
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_294
timestamp 1649977179
transform 1 0 28152 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_300
timestamp 1649977179
transform 1 0 28704 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_312
timestamp 1649977179
transform 1 0 29808 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_324
timestamp 1649977179
transform 1 0 30912 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_354
timestamp 1649977179
transform 1 0 33672 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_366
timestamp 1649977179
transform 1 0 34776 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_378
timestamp 1649977179
transform 1 0 35880 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1649977179
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_413
timestamp 1649977179
transform 1 0 39100 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_419
timestamp 1649977179
transform 1 0 39652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1649977179
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1649977179
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1649977179
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1649977179
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1649977179
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1649977179
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1649977179
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1649977179
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1649977179
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1649977179
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1649977179
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1649977179
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_565
timestamp 1649977179
transform 1 0 53084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_577
timestamp 1649977179
transform 1 0 54188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_589
timestamp 1649977179
transform 1 0 55292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_601
timestamp 1649977179
transform 1 0 56396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_613
timestamp 1649977179
transform 1 0 57500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_621
timestamp 1649977179
transform 1 0 58236 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_261
timestamp 1649977179
transform 1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_284
timestamp 1649977179
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_290
timestamp 1649977179
transform 1 0 27784 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1649977179
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_385
timestamp 1649977179
transform 1 0 36524 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_397
timestamp 1649977179
transform 1 0 37628 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_409
timestamp 1649977179
transform 1 0 38732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_417
timestamp 1649977179
transform 1 0 39468 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_441
timestamp 1649977179
transform 1 0 41676 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_453
timestamp 1649977179
transform 1 0 42780 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_465
timestamp 1649977179
transform 1 0 43884 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1649977179
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1649977179
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1649977179
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1649977179
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1649977179
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1649977179
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1649977179
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1649977179
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1649977179
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_265
timestamp 1649977179
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1649977179
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_284
timestamp 1649977179
transform 1 0 27232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_296
timestamp 1649977179
transform 1 0 28336 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_306
timestamp 1649977179
transform 1 0 29256 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_318
timestamp 1649977179
transform 1 0 30360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_322
timestamp 1649977179
transform 1 0 30728 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_330
timestamp 1649977179
transform 1 0 31464 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_363
timestamp 1649977179
transform 1 0 34500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1649977179
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_400
timestamp 1649977179
transform 1 0 37904 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_408
timestamp 1649977179
transform 1 0 38640 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_430
timestamp 1649977179
transform 1 0 40664 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_442
timestamp 1649977179
transform 1 0 41768 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_469
timestamp 1649977179
transform 1 0 44252 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_481
timestamp 1649977179
transform 1 0 45356 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_493
timestamp 1649977179
transform 1 0 46460 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_501
timestamp 1649977179
transform 1 0 47196 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_520
timestamp 1649977179
transform 1 0 48944 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_526
timestamp 1649977179
transform 1 0 49496 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_538
timestamp 1649977179
transform 1 0 50600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_550
timestamp 1649977179
transform 1 0 51704 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_558
timestamp 1649977179
transform 1 0 52440 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_260
timestamp 1649977179
transform 1 0 25024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_270
timestamp 1649977179
transform 1 0 25944 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_280
timestamp 1649977179
transform 1 0 26864 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1649977179
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_311
timestamp 1649977179
transform 1 0 29716 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_319
timestamp 1649977179
transform 1 0 30452 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_327
timestamp 1649977179
transform 1 0 31188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1649977179
transform 1 0 32108 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_353
timestamp 1649977179
transform 1 0 33580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_359
timestamp 1649977179
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_373
timestamp 1649977179
transform 1 0 35420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_385
timestamp 1649977179
transform 1 0 36524 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_393
timestamp 1649977179
transform 1 0 37260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_399
timestamp 1649977179
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_407
timestamp 1649977179
transform 1 0 38548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_424
timestamp 1649977179
transform 1 0 40112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_432
timestamp 1649977179
transform 1 0 40848 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_436
timestamp 1649977179
transform 1 0 41216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_440
timestamp 1649977179
transform 1 0 41584 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_461
timestamp 1649977179
transform 1 0 43516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_473
timestamp 1649977179
transform 1 0 44620 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_13
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_25
timestamp 1649977179
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_37
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1649977179
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_211
timestamp 1649977179
transform 1 0 20516 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_227
timestamp 1649977179
transform 1 0 21988 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_239
timestamp 1649977179
transform 1 0 23092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_251
timestamp 1649977179
transform 1 0 24196 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_259
timestamp 1649977179
transform 1 0 24932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_262
timestamp 1649977179
transform 1 0 25208 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_268
timestamp 1649977179
transform 1 0 25760 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp 1649977179
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_297
timestamp 1649977179
transform 1 0 28428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_319
timestamp 1649977179
transform 1 0 30452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_326
timestamp 1649977179
transform 1 0 31096 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1649977179
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_343
timestamp 1649977179
transform 1 0 32660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_370
timestamp 1649977179
transform 1 0 35144 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_378
timestamp 1649977179
transform 1 0 35880 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1649977179
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_400
timestamp 1649977179
transform 1 0 37904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_408
timestamp 1649977179
transform 1 0 38640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_432
timestamp 1649977179
transform 1 0 40848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1649977179
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_455
timestamp 1649977179
transform 1 0 42964 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_467
timestamp 1649977179
transform 1 0 44068 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_479
timestamp 1649977179
transform 1 0 45172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_491
timestamp 1649977179
transform 1 0 46276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_271
timestamp 1649977179
transform 1 0 26036 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_283
timestamp 1649977179
transform 1 0 27140 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_292
timestamp 1649977179
transform 1 0 27968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_296
timestamp 1649977179
transform 1 0 28336 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1649977179
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1649977179
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_331
timestamp 1649977179
transform 1 0 31556 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_339
timestamp 1649977179
transform 1 0 32292 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1649977179
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_430
timestamp 1649977179
transform 1 0 40664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_441
timestamp 1649977179
transform 1 0 41676 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_447
timestamp 1649977179
transform 1 0 42228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_454
timestamp 1649977179
transform 1 0 42872 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_463
timestamp 1649977179
transform 1 0 43700 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_471
timestamp 1649977179
transform 1 0 44436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_202
timestamp 1649977179
transform 1 0 19688 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_214
timestamp 1649977179
transform 1 0 20792 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1649977179
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_290
timestamp 1649977179
transform 1 0 27784 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_300
timestamp 1649977179
transform 1 0 28704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_308
timestamp 1649977179
transform 1 0 29440 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_314
timestamp 1649977179
transform 1 0 29992 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_322
timestamp 1649977179
transform 1 0 30728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_330
timestamp 1649977179
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_370
timestamp 1649977179
transform 1 0 35144 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_382
timestamp 1649977179
transform 1 0 36248 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1649977179
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_397
timestamp 1649977179
transform 1 0 37628 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_401
timestamp 1649977179
transform 1 0 37996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_416
timestamp 1649977179
transform 1 0 39376 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_420
timestamp 1649977179
transform 1 0 39744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_428
timestamp 1649977179
transform 1 0 40480 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_432
timestamp 1649977179
transform 1 0 40848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_437
timestamp 1649977179
transform 1 0 41308 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_444
timestamp 1649977179
transform 1 0 41952 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_458
timestamp 1649977179
transform 1 0 43240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_469
timestamp 1649977179
transform 1 0 44252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_475
timestamp 1649977179
transform 1 0 44804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_491
timestamp 1649977179
transform 1 0 46276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_201
timestamp 1649977179
transform 1 0 19596 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_210
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_225
timestamp 1649977179
transform 1 0 21804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_237
timestamp 1649977179
transform 1 0 22908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1649977179
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_288
timestamp 1649977179
transform 1 0 27600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_299
timestamp 1649977179
transform 1 0 28612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_312
timestamp 1649977179
transform 1 0 29808 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_318
timestamp 1649977179
transform 1 0 30360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_324
timestamp 1649977179
transform 1 0 30912 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_334
timestamp 1649977179
transform 1 0 31832 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_340
timestamp 1649977179
transform 1 0 32384 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_348
timestamp 1649977179
transform 1 0 33120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_354
timestamp 1649977179
transform 1 0 33672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1649977179
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_367
timestamp 1649977179
transform 1 0 34868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_371
timestamp 1649977179
transform 1 0 35236 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_392
timestamp 1649977179
transform 1 0 37168 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_400
timestamp 1649977179
transform 1 0 37904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_405
timestamp 1649977179
transform 1 0 38364 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_414
timestamp 1649977179
transform 1 0 39192 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_429
timestamp 1649977179
transform 1 0 40572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_435
timestamp 1649977179
transform 1 0 41124 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_441
timestamp 1649977179
transform 1 0 41676 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_454
timestamp 1649977179
transform 1 0 42872 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_466
timestamp 1649977179
transform 1 0 43976 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_474
timestamp 1649977179
transform 1 0 44712 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_479
timestamp 1649977179
transform 1 0 45172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_485
timestamp 1649977179
transform 1 0 45724 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_495
timestamp 1649977179
transform 1 0 46644 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_213
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_218
timestamp 1649977179
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_234
timestamp 1649977179
transform 1 0 22632 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_246
timestamp 1649977179
transform 1 0 23736 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_258
timestamp 1649977179
transform 1 0 24840 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1649977179
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1649977179
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_288
timestamp 1649977179
transform 1 0 27600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_299
timestamp 1649977179
transform 1 0 28612 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_308
timestamp 1649977179
transform 1 0 29440 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_315
timestamp 1649977179
transform 1 0 30084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp 1649977179
transform 1 0 30820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1649977179
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_344
timestamp 1649977179
transform 1 0 32752 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_356
timestamp 1649977179
transform 1 0 33856 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_367
timestamp 1649977179
transform 1 0 34868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_379
timestamp 1649977179
transform 1 0 35972 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1649977179
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_399
timestamp 1649977179
transform 1 0 37812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_424
timestamp 1649977179
transform 1 0 40112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_432
timestamp 1649977179
transform 1 0 40848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_439
timestamp 1649977179
transform 1 0 41492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_469
timestamp 1649977179
transform 1 0 44252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_476
timestamp 1649977179
transform 1 0 44896 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_484
timestamp 1649977179
transform 1 0 45632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_490
timestamp 1649977179
transform 1 0 46184 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_498
timestamp 1649977179
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_214
timestamp 1649977179
transform 1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_220
timestamp 1649977179
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_232
timestamp 1649977179
transform 1 0 22448 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1649977179
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_282
timestamp 1649977179
transform 1 0 27048 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_296
timestamp 1649977179
transform 1 0 28336 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1649977179
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_313
timestamp 1649977179
transform 1 0 29900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_324
timestamp 1649977179
transform 1 0 30912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_328
timestamp 1649977179
transform 1 0 31280 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_335
timestamp 1649977179
transform 1 0 31924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_353
timestamp 1649977179
transform 1 0 33580 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1649977179
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_386
timestamp 1649977179
transform 1 0 36616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_410
timestamp 1649977179
transform 1 0 38824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1649977179
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_444
timestamp 1649977179
transform 1 0 41952 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_468
timestamp 1649977179
transform 1 0 44160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_484
timestamp 1649977179
transform 1 0 45632 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_494
timestamp 1649977179
transform 1 0 46552 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_503
timestamp 1649977179
transform 1 0 47380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_515
timestamp 1649977179
transform 1 0 48484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_527
timestamp 1649977179
transform 1 0 49588 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_609
timestamp 1649977179
transform 1 0 57132 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_621
timestamp 1649977179
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_201
timestamp 1649977179
transform 1 0 19596 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_210
timestamp 1649977179
transform 1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_287
timestamp 1649977179
transform 1 0 27508 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_302
timestamp 1649977179
transform 1 0 28888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_309
timestamp 1649977179
transform 1 0 29532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_325
timestamp 1649977179
transform 1 0 31004 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1649977179
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_344
timestamp 1649977179
transform 1 0 32752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_350
timestamp 1649977179
transform 1 0 33304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_372
timestamp 1649977179
transform 1 0 35328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_378
timestamp 1649977179
transform 1 0 35880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1649977179
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_400
timestamp 1649977179
transform 1 0 37904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_411
timestamp 1649977179
transform 1 0 38916 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_426
timestamp 1649977179
transform 1 0 40296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_434
timestamp 1649977179
transform 1 0 41032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_451
timestamp 1649977179
transform 1 0 42596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_459
timestamp 1649977179
transform 1 0 43332 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_474
timestamp 1649977179
transform 1 0 44712 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_489
timestamp 1649977179
transform 1 0 46092 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_496
timestamp 1649977179
transform 1 0 46736 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_591
timestamp 1649977179
transform 1 0 55476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_603
timestamp 1649977179
transform 1 0 56580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_18
timestamp 1649977179
transform 1 0 2760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_167
timestamp 1649977179
transform 1 0 16468 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_201
timestamp 1649977179
transform 1 0 19596 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_211
timestamp 1649977179
transform 1 0 20516 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_217
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_223
timestamp 1649977179
transform 1 0 21620 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_235
timestamp 1649977179
transform 1 0 22724 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_247
timestamp 1649977179
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_269
timestamp 1649977179
transform 1 0 25852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_280
timestamp 1649977179
transform 1 0 26864 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_287
timestamp 1649977179
transform 1 0 27508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_298
timestamp 1649977179
transform 1 0 28520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_316
timestamp 1649977179
transform 1 0 30176 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_324
timestamp 1649977179
transform 1 0 30912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_332
timestamp 1649977179
transform 1 0 31648 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_360
timestamp 1649977179
transform 1 0 34224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_374
timestamp 1649977179
transform 1 0 35512 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1649977179
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_414
timestamp 1649977179
transform 1 0 39192 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_427
timestamp 1649977179
transform 1 0 40388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_435
timestamp 1649977179
transform 1 0 41124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_456
timestamp 1649977179
transform 1 0 43056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_460
timestamp 1649977179
transform 1 0 43424 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_464
timestamp 1649977179
transform 1 0 43792 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_472
timestamp 1649977179
transform 1 0 44528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_486
timestamp 1649977179
transform 1 0 45816 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_492
timestamp 1649977179
transform 1 0 46368 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_504
timestamp 1649977179
transform 1 0 47472 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_514
timestamp 1649977179
transform 1 0 48392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_526
timestamp 1649977179
transform 1 0 49496 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_537
timestamp 1649977179
transform 1 0 50508 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_543
timestamp 1649977179
transform 1 0 51060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_555
timestamp 1649977179
transform 1 0 52164 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_567
timestamp 1649977179
transform 1 0 53268 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_579
timestamp 1649977179
transform 1 0 54372 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_612
timestamp 1649977179
transform 1 0 57408 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_624
timestamp 1649977179
transform 1 0 58512 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1649977179
transform 1 0 18032 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1649977179
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_227
timestamp 1649977179
transform 1 0 21988 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_239
timestamp 1649977179
transform 1 0 23092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_272
timestamp 1649977179
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_302
timestamp 1649977179
transform 1 0 28888 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_310
timestamp 1649977179
transform 1 0 29624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1649977179
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_345
timestamp 1649977179
transform 1 0 32844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_353
timestamp 1649977179
transform 1 0 33580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_375
timestamp 1649977179
transform 1 0 35604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_383
timestamp 1649977179
transform 1 0 36340 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_397
timestamp 1649977179
transform 1 0 37628 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_425
timestamp 1649977179
transform 1 0 40204 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_434
timestamp 1649977179
transform 1 0 41032 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_442
timestamp 1649977179
transform 1 0 41768 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_456
timestamp 1649977179
transform 1 0 43056 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_462
timestamp 1649977179
transform 1 0 43608 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_470
timestamp 1649977179
transform 1 0 44344 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_475
timestamp 1649977179
transform 1 0 44804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_487
timestamp 1649977179
transform 1 0 45908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_499
timestamp 1649977179
transform 1 0 47012 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_512
timestamp 1649977179
transform 1 0 48208 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_518
timestamp 1649977179
transform 1 0 48760 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_539
timestamp 1649977179
transform 1 0 50692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_555
timestamp 1649977179
transform 1 0 52164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_577
timestamp 1649977179
transform 1 0 54188 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_598
timestamp 1649977179
transform 1 0 56120 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_610
timestamp 1649977179
transform 1 0 57224 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_621
timestamp 1649977179
transform 1 0 58236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_159
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_180
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_186
timestamp 1649977179
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1649977179
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_211
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_215
timestamp 1649977179
transform 1 0 20884 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_219
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_227
timestamp 1649977179
transform 1 0 21988 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1649977179
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_257
timestamp 1649977179
transform 1 0 24748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_279
timestamp 1649977179
transform 1 0 26772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_315
timestamp 1649977179
transform 1 0 30084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_323
timestamp 1649977179
transform 1 0 30820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_339
timestamp 1649977179
transform 1 0 32292 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_351
timestamp 1649977179
transform 1 0 33396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_355
timestamp 1649977179
transform 1 0 33764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1649977179
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_385
timestamp 1649977179
transform 1 0 36524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_409
timestamp 1649977179
transform 1 0 38732 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1649977179
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_430
timestamp 1649977179
transform 1 0 40664 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_438
timestamp 1649977179
transform 1 0 41400 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_459
timestamp 1649977179
transform 1 0 43332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_465
timestamp 1649977179
transform 1 0 43884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_471
timestamp 1649977179
transform 1 0 44436 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_485
timestamp 1649977179
transform 1 0 45724 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_497
timestamp 1649977179
transform 1 0 46828 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_509
timestamp 1649977179
transform 1 0 47932 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_515
timestamp 1649977179
transform 1 0 48484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_527
timestamp 1649977179
transform 1 0 49588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_541
timestamp 1649977179
transform 1 0 50876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_553
timestamp 1649977179
transform 1 0 51980 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_563
timestamp 1649977179
transform 1 0 52900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_575
timestamp 1649977179
transform 1 0 54004 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_593
timestamp 1649977179
transform 1 0 55660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_596
timestamp 1649977179
transform 1 0 55936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_620
timestamp 1649977179
transform 1 0 58144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_624
timestamp 1649977179
transform 1 0 58512 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1649977179
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_175
timestamp 1649977179
transform 1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_187
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_190
timestamp 1649977179
transform 1 0 18584 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_214
timestamp 1649977179
transform 1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1649977179
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_230
timestamp 1649977179
transform 1 0 22264 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_236
timestamp 1649977179
transform 1 0 22816 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_258
timestamp 1649977179
transform 1 0 24840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_262
timestamp 1649977179
transform 1 0 25208 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1649977179
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_302
timestamp 1649977179
transform 1 0 28888 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_308
timestamp 1649977179
transform 1 0 29440 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1649977179
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_344
timestamp 1649977179
transform 1 0 32752 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_352
timestamp 1649977179
transform 1 0 33488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_375
timestamp 1649977179
transform 1 0 35604 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_386
timestamp 1649977179
transform 1 0 36616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_400
timestamp 1649977179
transform 1 0 37904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_408
timestamp 1649977179
transform 1 0 38640 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_432
timestamp 1649977179
transform 1 0 40848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_440
timestamp 1649977179
transform 1 0 41584 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_453
timestamp 1649977179
transform 1 0 42780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_465
timestamp 1649977179
transform 1 0 43884 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_476
timestamp 1649977179
transform 1 0 44896 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_482
timestamp 1649977179
transform 1 0 45448 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_494
timestamp 1649977179
transform 1 0 46552 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_502
timestamp 1649977179
transform 1 0 47288 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_508
timestamp 1649977179
transform 1 0 47840 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_514
timestamp 1649977179
transform 1 0 48392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_521
timestamp 1649977179
transform 1 0 49036 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_554
timestamp 1649977179
transform 1 0 52072 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_569
timestamp 1649977179
transform 1 0 53452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_581
timestamp 1649977179
transform 1 0 54556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_593
timestamp 1649977179
transform 1 0 55660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_605
timestamp 1649977179
transform 1 0 56764 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_613
timestamp 1649977179
transform 1 0 57500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_117
timestamp 1649977179
transform 1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_123
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_129
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_143
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1649977179
transform 1 0 15364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_179
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_200
timestamp 1649977179
transform 1 0 19504 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1649977179
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_256
timestamp 1649977179
transform 1 0 24656 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_262
timestamp 1649977179
transform 1 0 25208 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_276
timestamp 1649977179
transform 1 0 26496 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_282
timestamp 1649977179
transform 1 0 27048 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_290
timestamp 1649977179
transform 1 0 27784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_294
timestamp 1649977179
transform 1 0 28152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_316
timestamp 1649977179
transform 1 0 30176 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_325
timestamp 1649977179
transform 1 0 31004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_347
timestamp 1649977179
transform 1 0 33028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_353
timestamp 1649977179
transform 1 0 33580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_359
timestamp 1649977179
transform 1 0 34132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_395
timestamp 1649977179
transform 1 0 37444 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1649977179
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_414
timestamp 1649977179
transform 1 0 39192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_429
timestamp 1649977179
transform 1 0 40572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_453
timestamp 1649977179
transform 1 0 42780 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_463
timestamp 1649977179
transform 1 0 43700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_484
timestamp 1649977179
transform 1 0 45632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_496
timestamp 1649977179
transform 1 0 46736 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_500
timestamp 1649977179
transform 1 0 47104 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_504
timestamp 1649977179
transform 1 0 47472 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_514
timestamp 1649977179
transform 1 0 48392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_518
timestamp 1649977179
transform 1 0 48760 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_526
timestamp 1649977179
transform 1 0 49496 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_553
timestamp 1649977179
transform 1 0 51980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_561
timestamp 1649977179
transform 1 0 52716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_568
timestamp 1649977179
transform 1 0 53360 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_575
timestamp 1649977179
transform 1 0 54004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_621
timestamp 1649977179
transform 1 0 58236 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_128
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_134
timestamp 1649977179
transform 1 0 13432 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_173
timestamp 1649977179
transform 1 0 17020 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_183
timestamp 1649977179
transform 1 0 17940 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_239
timestamp 1649977179
transform 1 0 23092 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_263
timestamp 1649977179
transform 1 0 25300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_269
timestamp 1649977179
transform 1 0 25852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1649977179
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_314
timestamp 1649977179
transform 1 0 29992 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_325
timestamp 1649977179
transform 1 0 31004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1649977179
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_343
timestamp 1649977179
transform 1 0 32660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_357
timestamp 1649977179
transform 1 0 33948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_368
timestamp 1649977179
transform 1 0 34960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_377
timestamp 1649977179
transform 1 0 35788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_381
timestamp 1649977179
transform 1 0 36156 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_414
timestamp 1649977179
transform 1 0 39192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_425
timestamp 1649977179
transform 1 0 40204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_432
timestamp 1649977179
transform 1 0 40848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1649977179
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_452
timestamp 1649977179
transform 1 0 42688 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_460
timestamp 1649977179
transform 1 0 43424 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_465
timestamp 1649977179
transform 1 0 43884 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_492
timestamp 1649977179
transform 1 0 46368 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_514
timestamp 1649977179
transform 1 0 48392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_523
timestamp 1649977179
transform 1 0 49220 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_531
timestamp 1649977179
transform 1 0 49956 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_536
timestamp 1649977179
transform 1 0 50416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_550
timestamp 1649977179
transform 1 0 51704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_556
timestamp 1649977179
transform 1 0 52256 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_570
timestamp 1649977179
transform 1 0 53544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_578
timestamp 1649977179
transform 1 0 54280 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_582
timestamp 1649977179
transform 1 0 54648 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_590
timestamp 1649977179
transform 1 0 55384 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_596
timestamp 1649977179
transform 1 0 55936 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_604
timestamp 1649977179
transform 1 0 56672 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_167
timestamp 1649977179
transform 1 0 16468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1649977179
transform 1 0 20424 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1649977179
transform 1 0 22632 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1649977179
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1649977179
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_273
timestamp 1649977179
transform 1 0 26220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1649977179
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_313
timestamp 1649977179
transform 1 0 29900 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_320
timestamp 1649977179
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_324
timestamp 1649977179
transform 1 0 30912 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_331
timestamp 1649977179
transform 1 0 31556 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_351
timestamp 1649977179
transform 1 0 33396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1649977179
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_368
timestamp 1649977179
transform 1 0 34960 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_372
timestamp 1649977179
transform 1 0 35328 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_383
timestamp 1649977179
transform 1 0 36340 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_391
timestamp 1649977179
transform 1 0 37076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_399
timestamp 1649977179
transform 1 0 37812 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_410
timestamp 1649977179
transform 1 0 38824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1649977179
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_427
timestamp 1649977179
transform 1 0 40388 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_447
timestamp 1649977179
transform 1 0 42228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_455
timestamp 1649977179
transform 1 0 42964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_463
timestamp 1649977179
transform 1 0 43700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_472
timestamp 1649977179
transform 1 0 44528 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_497
timestamp 1649977179
transform 1 0 46828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_521
timestamp 1649977179
transform 1 0 49036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_528
timestamp 1649977179
transform 1 0 49680 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_546
timestamp 1649977179
transform 1 0 51336 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_570
timestamp 1649977179
transform 1 0 53544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_580
timestamp 1649977179
transform 1 0 54464 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_609
timestamp 1649977179
transform 1 0 57132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_621
timestamp 1649977179
transform 1 0 58236 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_76
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_126
timestamp 1649977179
transform 1 0 12696 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_132
timestamp 1649977179
transform 1 0 13248 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1649977179
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_173
timestamp 1649977179
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_195
timestamp 1649977179
transform 1 0 19044 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_216
timestamp 1649977179
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_248
timestamp 1649977179
transform 1 0 23920 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1649977179
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_283
timestamp 1649977179
transform 1 0 27140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_290
timestamp 1649977179
transform 1 0 27784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_315
timestamp 1649977179
transform 1 0 30084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_328
timestamp 1649977179
transform 1 0 31280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_344
timestamp 1649977179
transform 1 0 32752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_350
timestamp 1649977179
transform 1 0 33304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_354
timestamp 1649977179
transform 1 0 33672 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_375
timestamp 1649977179
transform 1 0 35604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_384
timestamp 1649977179
transform 1 0 36432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_414
timestamp 1649977179
transform 1 0 39192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_420
timestamp 1649977179
transform 1 0 39744 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_426
timestamp 1649977179
transform 1 0 40296 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_444
timestamp 1649977179
transform 1 0 41952 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_452
timestamp 1649977179
transform 1 0 42688 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_464
timestamp 1649977179
transform 1 0 43792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_470
timestamp 1649977179
transform 1 0 44344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_477
timestamp 1649977179
transform 1 0 44988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_493
timestamp 1649977179
transform 1 0 46460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_500
timestamp 1649977179
transform 1 0 47104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_507
timestamp 1649977179
transform 1 0 47748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_518
timestamp 1649977179
transform 1 0 48760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_526
timestamp 1649977179
transform 1 0 49496 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_555
timestamp 1649977179
transform 1 0 52164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_569
timestamp 1649977179
transform 1 0 53452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_593
timestamp 1649977179
transform 1 0 55660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_601
timestamp 1649977179
transform 1 0 56396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_612
timestamp 1649977179
transform 1 0 57408 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_621
timestamp 1649977179
transform 1 0 58236 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_73
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1649977179
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1649977179
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1649977179
transform 1 0 16100 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_200
timestamp 1649977179
transform 1 0 19504 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_224
timestamp 1649977179
transform 1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1649977179
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_256
timestamp 1649977179
transform 1 0 24656 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1649977179
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_291
timestamp 1649977179
transform 1 0 27876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1649977179
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_312
timestamp 1649977179
transform 1 0 29808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_316
timestamp 1649977179
transform 1 0 30176 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_346
timestamp 1649977179
transform 1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_352
timestamp 1649977179
transform 1 0 33488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_358
timestamp 1649977179
transform 1 0 34040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_371
timestamp 1649977179
transform 1 0 35236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_396
timestamp 1649977179
transform 1 0 37536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_403
timestamp 1649977179
transform 1 0 38180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_411
timestamp 1649977179
transform 1 0 38916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1649977179
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_425
timestamp 1649977179
transform 1 0 40204 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_429
timestamp 1649977179
transform 1 0 40572 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_447
timestamp 1649977179
transform 1 0 42228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_465
timestamp 1649977179
transform 1 0 43884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_472
timestamp 1649977179
transform 1 0 44528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_485
timestamp 1649977179
transform 1 0 45724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_492
timestamp 1649977179
transform 1 0 46368 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_498
timestamp 1649977179
transform 1 0 46920 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_505
timestamp 1649977179
transform 1 0 47564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_509
timestamp 1649977179
transform 1 0 47932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_514
timestamp 1649977179
transform 1 0 48392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_524
timestamp 1649977179
transform 1 0 49312 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_536
timestamp 1649977179
transform 1 0 50416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_543
timestamp 1649977179
transform 1 0 51060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_575
timestamp 1649977179
transform 1 0 54004 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_583
timestamp 1649977179
transform 1 0 54740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_621
timestamp 1649977179
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_64
timestamp 1649977179
transform 1 0 6992 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_70
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_84
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1649977179
transform 1 0 11868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1649977179
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_131
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_143
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_171
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1649977179
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_209
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_284
timestamp 1649977179
transform 1 0 27232 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_310
timestamp 1649977179
transform 1 0 29624 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_316
timestamp 1649977179
transform 1 0 30176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_321
timestamp 1649977179
transform 1 0 30636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1649977179
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_350
timestamp 1649977179
transform 1 0 33304 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_377
timestamp 1649977179
transform 1 0 35788 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_389
timestamp 1649977179
transform 1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_426
timestamp 1649977179
transform 1 0 40296 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_444
timestamp 1649977179
transform 1 0 41952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_463
timestamp 1649977179
transform 1 0 43700 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_470
timestamp 1649977179
transform 1 0 44344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_474
timestamp 1649977179
transform 1 0 44712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_482
timestamp 1649977179
transform 1 0 45448 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_490
timestamp 1649977179
transform 1 0 46184 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_525
timestamp 1649977179
transform 1 0 49404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_533
timestamp 1649977179
transform 1 0 50140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_540
timestamp 1649977179
transform 1 0 50784 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_556
timestamp 1649977179
transform 1 0 52256 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_569
timestamp 1649977179
transform 1 0 53452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_576
timestamp 1649977179
transform 1 0 54096 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_583
timestamp 1649977179
transform 1 0 54740 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_595
timestamp 1649977179
transform 1 0 55844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_604
timestamp 1649977179
transform 1 0 56672 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_612
timestamp 1649977179
transform 1 0 57408 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_620
timestamp 1649977179
transform 1 0 58144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_624
timestamp 1649977179
transform 1 0 58512 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_49
timestamp 1649977179
transform 1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_54
timestamp 1649977179
transform 1 0 6072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_61
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_73
timestamp 1649977179
transform 1 0 7820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_90
timestamp 1649977179
transform 1 0 9384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_125
timestamp 1649977179
transform 1 0 12604 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_129
timestamp 1649977179
transform 1 0 12972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1649977179
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_203
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_207
timestamp 1649977179
transform 1 0 20148 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_211
timestamp 1649977179
transform 1 0 20516 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_222
timestamp 1649977179
transform 1 0 21528 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1649977179
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_273
timestamp 1649977179
transform 1 0 26220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1649977179
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_284
timestamp 1649977179
transform 1 0 27232 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1649977179
transform 1 0 28520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1649977179
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_316
timestamp 1649977179
transform 1 0 30176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_340
timestamp 1649977179
transform 1 0 32384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_346
timestamp 1649977179
transform 1 0 32936 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_354
timestamp 1649977179
transform 1 0 33672 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_369
timestamp 1649977179
transform 1 0 35052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_390
timestamp 1649977179
transform 1 0 36984 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_394
timestamp 1649977179
transform 1 0 37352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_397
timestamp 1649977179
transform 1 0 37628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_414
timestamp 1649977179
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_425
timestamp 1649977179
transform 1 0 40204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_429
timestamp 1649977179
transform 1 0 40572 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_447
timestamp 1649977179
transform 1 0 42228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_465
timestamp 1649977179
transform 1 0 43884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_472
timestamp 1649977179
transform 1 0 44528 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_483
timestamp 1649977179
transform 1 0 45540 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_491
timestamp 1649977179
transform 1 0 46276 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_502
timestamp 1649977179
transform 1 0 47288 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_516
timestamp 1649977179
transform 1 0 48576 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_523
timestamp 1649977179
transform 1 0 49220 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_544
timestamp 1649977179
transform 1 0 51152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_555
timestamp 1649977179
transform 1 0 52164 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_563
timestamp 1649977179
transform 1 0 52900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_571
timestamp 1649977179
transform 1 0 53636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_579
timestamp 1649977179
transform 1 0 54372 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1649977179
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_46
timestamp 1649977179
transform 1 0 5336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_63
timestamp 1649977179
transform 1 0 6900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_70
timestamp 1649977179
transform 1 0 7544 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_84
timestamp 1649977179
transform 1 0 8832 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_116
timestamp 1649977179
transform 1 0 11776 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_173
timestamp 1649977179
transform 1 0 17020 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_198
timestamp 1649977179
transform 1 0 19320 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_206
timestamp 1649977179
transform 1 0 20056 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1649977179
transform 1 0 23644 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_252
timestamp 1649977179
transform 1 0 24288 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1649977179
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_288
timestamp 1649977179
transform 1 0 27600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_295
timestamp 1649977179
transform 1 0 28244 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_301
timestamp 1649977179
transform 1 0 28796 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_323
timestamp 1649977179
transform 1 0 30820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_340
timestamp 1649977179
transform 1 0 32384 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_346
timestamp 1649977179
transform 1 0 32936 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_352
timestamp 1649977179
transform 1 0 33488 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1649977179
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_381
timestamp 1649977179
transform 1 0 36156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1649977179
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_413
timestamp 1649977179
transform 1 0 39100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_420
timestamp 1649977179
transform 1 0 39744 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_426
timestamp 1649977179
transform 1 0 40296 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_444
timestamp 1649977179
transform 1 0 41952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_453
timestamp 1649977179
transform 1 0 42780 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_459
timestamp 1649977179
transform 1 0 43332 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_481
timestamp 1649977179
transform 1 0 45356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_498
timestamp 1649977179
transform 1 0 46920 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_511
timestamp 1649977179
transform 1 0 48116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_519
timestamp 1649977179
transform 1 0 48852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_540
timestamp 1649977179
transform 1 0 50784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_551
timestamp 1649977179
transform 1 0 51796 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_567
timestamp 1649977179
transform 1 0 53268 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_575
timestamp 1649977179
transform 1 0 54004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_583
timestamp 1649977179
transform 1 0 54740 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_607
timestamp 1649977179
transform 1 0 56948 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_54
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_71
timestamp 1649977179
transform 1 0 7636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_89
timestamp 1649977179
transform 1 0 9292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_96
timestamp 1649977179
transform 1 0 9936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1649977179
transform 1 0 10304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1649977179
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_132
timestamp 1649977179
transform 1 0 13248 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_148
timestamp 1649977179
transform 1 0 14720 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_173
timestamp 1649977179
transform 1 0 17020 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_181
timestamp 1649977179
transform 1 0 17756 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1649977179
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1649977179
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_230
timestamp 1649977179
transform 1 0 22264 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1649977179
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_241
timestamp 1649977179
transform 1 0 23276 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1649977179
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_256
timestamp 1649977179
transform 1 0 24656 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_262
timestamp 1649977179
transform 1 0 25208 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_266
timestamp 1649977179
transform 1 0 25576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_290
timestamp 1649977179
transform 1 0 27784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_297
timestamp 1649977179
transform 1 0 28428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1649977179
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_330
timestamp 1649977179
transform 1 0 31464 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_338
timestamp 1649977179
transform 1 0 32200 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_351
timestamp 1649977179
transform 1 0 33396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1649977179
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_385
timestamp 1649977179
transform 1 0 36524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_392
timestamp 1649977179
transform 1 0 37168 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_400
timestamp 1649977179
transform 1 0 37904 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_408
timestamp 1649977179
transform 1 0 38640 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1649977179
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_428
timestamp 1649977179
transform 1 0 40480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_435
timestamp 1649977179
transform 1 0 41124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_439
timestamp 1649977179
transform 1 0 41492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_460
timestamp 1649977179
transform 1 0 43424 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_464
timestamp 1649977179
transform 1 0 43792 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_472
timestamp 1649977179
transform 1 0 44528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_498
timestamp 1649977179
transform 1 0 46920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_502
timestamp 1649977179
transform 1 0 47288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_507
timestamp 1649977179
transform 1 0 47748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_518
timestamp 1649977179
transform 1 0 48760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_526
timestamp 1649977179
transform 1 0 49496 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_536
timestamp 1649977179
transform 1 0 50416 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_542
timestamp 1649977179
transform 1 0 50968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_546
timestamp 1649977179
transform 1 0 51336 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_556
timestamp 1649977179
transform 1 0 52256 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_567
timestamp 1649977179
transform 1 0 53268 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_573
timestamp 1649977179
transform 1 0 53820 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_578
timestamp 1649977179
transform 1 0 54280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_584
timestamp 1649977179
transform 1 0 54832 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_597
timestamp 1649977179
transform 1 0 56028 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_620
timestamp 1649977179
transform 1 0 58144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_624
timestamp 1649977179
transform 1 0 58512 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_23
timestamp 1649977179
transform 1 0 3220 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1649977179
transform 1 0 3496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_32
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_60
timestamp 1649977179
transform 1 0 6624 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1649977179
transform 1 0 8832 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 1649977179
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_138
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_173
timestamp 1649977179
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_195
timestamp 1649977179
transform 1 0 19044 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_220
timestamp 1649977179
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_233
timestamp 1649977179
transform 1 0 22540 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_258
timestamp 1649977179
transform 1 0 24840 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1649977179
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_298
timestamp 1649977179
transform 1 0 28520 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1649977179
transform 1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_319
timestamp 1649977179
transform 1 0 30452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_323
timestamp 1649977179
transform 1 0 30820 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1649977179
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_357
timestamp 1649977179
transform 1 0 33948 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_365
timestamp 1649977179
transform 1 0 34684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_370
timestamp 1649977179
transform 1 0 35144 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_376
timestamp 1649977179
transform 1 0 35696 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1649977179
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_400
timestamp 1649977179
transform 1 0 37904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_404
timestamp 1649977179
transform 1 0 38272 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_408
timestamp 1649977179
transform 1 0 38640 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_415
timestamp 1649977179
transform 1 0 39284 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_422
timestamp 1649977179
transform 1 0 39928 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_430
timestamp 1649977179
transform 1 0 40664 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_444
timestamp 1649977179
transform 1 0 41952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_469
timestamp 1649977179
transform 1 0 44252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_479
timestamp 1649977179
transform 1 0 45172 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_515
timestamp 1649977179
transform 1 0 48484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_524
timestamp 1649977179
transform 1 0 49312 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_530
timestamp 1649977179
transform 1 0 49864 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_536
timestamp 1649977179
transform 1 0 50416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_543
timestamp 1649977179
transform 1 0 51060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_556
timestamp 1649977179
transform 1 0 52256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_565
timestamp 1649977179
transform 1 0 53084 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_576
timestamp 1649977179
transform 1 0 54096 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_588
timestamp 1649977179
transform 1 0 55200 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_612
timestamp 1649977179
transform 1 0 57408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_21
timestamp 1649977179
transform 1 0 3036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_39
timestamp 1649977179
transform 1 0 4692 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_46
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_63
timestamp 1649977179
transform 1 0 6900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_98
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_107
timestamp 1649977179
transform 1 0 10948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_132
timestamp 1649977179
transform 1 0 13248 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1649977179
transform 1 0 14352 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_151
timestamp 1649977179
transform 1 0 14996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_158
timestamp 1649977179
transform 1 0 15640 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1649977179
transform 1 0 17940 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1649977179
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_218
timestamp 1649977179
transform 1 0 21160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_224
timestamp 1649977179
transform 1 0 21712 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1649977179
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_273
timestamp 1649977179
transform 1 0 26220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_280
timestamp 1649977179
transform 1 0 26864 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_284
timestamp 1649977179
transform 1 0 27232 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1649977179
transform 1 0 27600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_296
timestamp 1649977179
transform 1 0 28336 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1649977179
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_316
timestamp 1649977179
transform 1 0 30176 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_324
timestamp 1649977179
transform 1 0 30912 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1649977179
transform 1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1649977179
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_368
timestamp 1649977179
transform 1 0 34960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_375
timestamp 1649977179
transform 1 0 35604 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1649977179
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_410
timestamp 1649977179
transform 1 0 38824 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1649977179
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_425
timestamp 1649977179
transform 1 0 40204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_432
timestamp 1649977179
transform 1 0 40848 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_459
timestamp 1649977179
transform 1 0 43332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_467
timestamp 1649977179
transform 1 0 44068 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_509
timestamp 1649977179
transform 1 0 47932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_516
timestamp 1649977179
transform 1 0 48576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_540
timestamp 1649977179
transform 1 0 50784 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_546
timestamp 1649977179
transform 1 0 51336 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_568
timestamp 1649977179
transform 1 0 53360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_572
timestamp 1649977179
transform 1 0 53728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_579
timestamp 1649977179
transform 1 0 54372 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_596
timestamp 1649977179
transform 1 0 55936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_600
timestamp 1649977179
transform 1 0 56304 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1649977179
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_35
timestamp 1649977179
transform 1 0 4324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1649977179
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_64
timestamp 1649977179
transform 1 0 6992 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_72
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_101
timestamp 1649977179
transform 1 0 10396 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1649977179
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_136
timestamp 1649977179
transform 1 0 13616 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1649977179
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_190
timestamp 1649977179
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1649977179
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_228
timestamp 1649977179
transform 1 0 22080 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_262
timestamp 1649977179
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_269
timestamp 1649977179
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1649977179
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_283
timestamp 1649977179
transform 1 0 27140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_289
timestamp 1649977179
transform 1 0 27692 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_306
timestamp 1649977179
transform 1 0 29256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_323
timestamp 1649977179
transform 1 0 30820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1649977179
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_358
timestamp 1649977179
transform 1 0 34040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1649977179
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1649977179
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_413
timestamp 1649977179
transform 1 0 39100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_437
timestamp 1649977179
transform 1 0 41308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_444
timestamp 1649977179
transform 1 0 41952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_470
timestamp 1649977179
transform 1 0 44344 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_478
timestamp 1649977179
transform 1 0 45080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1649977179
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_512
timestamp 1649977179
transform 1 0 48208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_518
timestamp 1649977179
transform 1 0 48760 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_524
timestamp 1649977179
transform 1 0 49312 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_545
timestamp 1649977179
transform 1 0 51244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_549
timestamp 1649977179
transform 1 0 51612 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_556
timestamp 1649977179
transform 1 0 52256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_582
timestamp 1649977179
transform 1 0 54648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_592
timestamp 1649977179
transform 1 0 55568 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_598
timestamp 1649977179
transform 1 0 56120 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_612
timestamp 1649977179
transform 1 0 57408 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_620
timestamp 1649977179
transform 1 0 58144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_624
timestamp 1649977179
transform 1 0 58512 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_14
timestamp 1649977179
transform 1 0 2392 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1649977179
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_51
timestamp 1649977179
transform 1 0 5796 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1649977179
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1649977179
transform 1 0 9200 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1649977179
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1649977179
transform 1 0 14352 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_150
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_182
timestamp 1649977179
transform 1 0 17848 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_188
timestamp 1649977179
transform 1 0 18400 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1649977179
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_231
timestamp 1649977179
transform 1 0 22356 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_238
timestamp 1649977179
transform 1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_255
timestamp 1649977179
transform 1 0 24564 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_279
timestamp 1649977179
transform 1 0 26772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_287
timestamp 1649977179
transform 1 0 27508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1649977179
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_311
timestamp 1649977179
transform 1 0 29716 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_323
timestamp 1649977179
transform 1 0 30820 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_329
timestamp 1649977179
transform 1 0 31372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_354
timestamp 1649977179
transform 1 0 33672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1649977179
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_369
timestamp 1649977179
transform 1 0 35052 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_374
timestamp 1649977179
transform 1 0 35512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_398
timestamp 1649977179
transform 1 0 37720 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_405
timestamp 1649977179
transform 1 0 38364 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_411
timestamp 1649977179
transform 1 0 38916 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_416
timestamp 1649977179
transform 1 0 39376 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_434
timestamp 1649977179
transform 1 0 41032 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_441
timestamp 1649977179
transform 1 0 41676 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_447
timestamp 1649977179
transform 1 0 42228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_498
timestamp 1649977179
transform 1 0 46920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_509
timestamp 1649977179
transform 1 0 47932 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_523
timestamp 1649977179
transform 1 0 49220 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_540
timestamp 1649977179
transform 1 0 50784 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_548
timestamp 1649977179
transform 1 0 51520 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_552
timestamp 1649977179
transform 1 0 51888 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_559
timestamp 1649977179
transform 1 0 52532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_570
timestamp 1649977179
transform 1 0 53544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_580
timestamp 1649977179
transform 1 0 54464 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_597
timestamp 1649977179
transform 1 0 56028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_621
timestamp 1649977179
transform 1 0 58236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_20
timestamp 1649977179
transform 1 0 2944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_35
timestamp 1649977179
transform 1 0 4324 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_41
timestamp 1649977179
transform 1 0 4876 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_45
timestamp 1649977179
transform 1 0 5244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1649977179
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_60
timestamp 1649977179
transform 1 0 6624 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_84
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_116
timestamp 1649977179
transform 1 0 11776 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_142
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_155
timestamp 1649977179
transform 1 0 15364 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1649977179
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_190
timestamp 1649977179
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_214
timestamp 1649977179
transform 1 0 20792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1649977179
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1649977179
transform 1 0 27416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_299
timestamp 1649977179
transform 1 0 28612 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_310
timestamp 1649977179
transform 1 0 29624 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_325
timestamp 1649977179
transform 1 0 31004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1649977179
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_344
timestamp 1649977179
transform 1 0 32752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_352
timestamp 1649977179
transform 1 0 33488 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_358
timestamp 1649977179
transform 1 0 34040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_383
timestamp 1649977179
transform 1 0 36340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1649977179
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_407
timestamp 1649977179
transform 1 0 38548 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_436
timestamp 1649977179
transform 1 0 41216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_443
timestamp 1649977179
transform 1 0 41860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_463
timestamp 1649977179
transform 1 0 43700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_474
timestamp 1649977179
transform 1 0 44712 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_478
timestamp 1649977179
transform 1 0 45080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_500
timestamp 1649977179
transform 1 0 47104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_513
timestamp 1649977179
transform 1 0 48300 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_519
timestamp 1649977179
transform 1 0 48852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_548
timestamp 1649977179
transform 1 0 51520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_552
timestamp 1649977179
transform 1 0 51888 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_556
timestamp 1649977179
transform 1 0 52256 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_568
timestamp 1649977179
transform 1 0 53360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_574
timestamp 1649977179
transform 1 0 53912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_588
timestamp 1649977179
transform 1 0 55200 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_596
timestamp 1649977179
transform 1 0 55936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_605
timestamp 1649977179
transform 1 0 56764 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_613
timestamp 1649977179
transform 1 0 57500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_621
timestamp 1649977179
transform 1 0 58236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_16
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1649977179
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_42
timestamp 1649977179
transform 1 0 4968 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_94
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_101
timestamp 1649977179
transform 1 0 10396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_108
timestamp 1649977179
transform 1 0 11040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_154
timestamp 1649977179
transform 1 0 15272 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_183
timestamp 1649977179
transform 1 0 17940 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1649977179
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1649977179
transform 1 0 20424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_229
timestamp 1649977179
transform 1 0 22172 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_237
timestamp 1649977179
transform 1 0 22908 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1649977179
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_263
timestamp 1649977179
transform 1 0 25300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_280
timestamp 1649977179
transform 1 0 26864 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1649977179
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_331
timestamp 1649977179
transform 1 0 31556 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1649977179
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_388
timestamp 1649977179
transform 1 0 36800 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_405
timestamp 1649977179
transform 1 0 38364 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_441
timestamp 1649977179
transform 1 0 41676 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_447
timestamp 1649977179
transform 1 0 42228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_452
timestamp 1649977179
transform 1 0 42688 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1649977179
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_482
timestamp 1649977179
transform 1 0 45448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_507
timestamp 1649977179
transform 1 0 47748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_518
timestamp 1649977179
transform 1 0 48760 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_527
timestamp 1649977179
transform 1 0 49588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_536
timestamp 1649977179
transform 1 0 50416 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_542
timestamp 1649977179
transform 1 0 50968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_548
timestamp 1649977179
transform 1 0 51520 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_567
timestamp 1649977179
transform 1 0 53268 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_573
timestamp 1649977179
transform 1 0 53820 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_584
timestamp 1649977179
transform 1 0 54832 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_618
timestamp 1649977179
transform 1 0 57960 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_624
timestamp 1649977179
transform 1 0 58512 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_16
timestamp 1649977179
transform 1 0 2576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_22
timestamp 1649977179
transform 1 0 3128 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_46
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1649977179
transform 1 0 6808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_97
timestamp 1649977179
transform 1 0 10028 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_101
timestamp 1649977179
transform 1 0 10396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1649977179
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_155
timestamp 1649977179
transform 1 0 15364 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1649977179
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_171
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1649977179
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1649977179
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_196
timestamp 1649977179
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_199
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_210
timestamp 1649977179
transform 1 0 20424 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_228
timestamp 1649977179
transform 1 0 22080 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_252
timestamp 1649977179
transform 1 0 24288 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_259
timestamp 1649977179
transform 1 0 24932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1649977179
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1649977179
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 1649977179
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_309
timestamp 1649977179
transform 1 0 29532 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_320
timestamp 1649977179
transform 1 0 30544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_327
timestamp 1649977179
transform 1 0 31188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_357
timestamp 1649977179
transform 1 0 33948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1649977179
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_388
timestamp 1649977179
transform 1 0 36800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_406
timestamp 1649977179
transform 1 0 38456 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_434
timestamp 1649977179
transform 1 0 41032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_442
timestamp 1649977179
transform 1 0 41768 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_452
timestamp 1649977179
transform 1 0 42688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_459
timestamp 1649977179
transform 1 0 43332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_477
timestamp 1649977179
transform 1 0 44988 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_495
timestamp 1649977179
transform 1 0 46644 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_512
timestamp 1649977179
transform 1 0 48208 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_520
timestamp 1649977179
transform 1 0 48944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_545
timestamp 1649977179
transform 1 0 51244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_552
timestamp 1649977179
transform 1 0 51888 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_567
timestamp 1649977179
transform 1 0 53268 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_574
timestamp 1649977179
transform 1 0 53912 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_598
timestamp 1649977179
transform 1 0 56120 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_610
timestamp 1649977179
transform 1 0 57224 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1649977179
transform 1 0 2576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1649977179
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1649977179
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_92
timestamp 1649977179
transform 1 0 9568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1649977179
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1649977179
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_130
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_151
timestamp 1649977179
transform 1 0 14996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_155
timestamp 1649977179
transform 1 0 15364 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_169
timestamp 1649977179
transform 1 0 16652 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_186
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_205
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_212
timestamp 1649977179
transform 1 0 20608 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1649977179
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_228
timestamp 1649977179
transform 1 0 22080 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_236
timestamp 1649977179
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_242
timestamp 1649977179
transform 1 0 23368 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1649977179
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_261
timestamp 1649977179
transform 1 0 25116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_269
timestamp 1649977179
transform 1 0 25852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1649977179
transform 1 0 27416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_296
timestamp 1649977179
transform 1 0 28336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_300
timestamp 1649977179
transform 1 0 28704 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1649977179
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_312
timestamp 1649977179
transform 1 0 29808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_320
timestamp 1649977179
transform 1 0 30544 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_341
timestamp 1649977179
transform 1 0 32476 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_348
timestamp 1649977179
transform 1 0 33120 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_355
timestamp 1649977179
transform 1 0 33764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_381
timestamp 1649977179
transform 1 0 36156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 1649977179
transform 1 0 38088 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_410
timestamp 1649977179
transform 1 0 38824 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1649977179
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_441
timestamp 1649977179
transform 1 0 41676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_448
timestamp 1649977179
transform 1 0 42320 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_454
timestamp 1649977179
transform 1 0 42872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1649977179
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_491
timestamp 1649977179
transform 1 0 46276 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_499
timestamp 1649977179
transform 1 0 47012 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_521
timestamp 1649977179
transform 1 0 49036 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_528
timestamp 1649977179
transform 1 0 49680 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_539
timestamp 1649977179
transform 1 0 50692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_546
timestamp 1649977179
transform 1 0 51336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_568
timestamp 1649977179
transform 1 0 53360 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_576
timestamp 1649977179
transform 1 0 54096 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_596
timestamp 1649977179
transform 1 0 55936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_620
timestamp 1649977179
transform 1 0 58144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_624
timestamp 1649977179
transform 1 0 58512 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_14
timestamp 1649977179
transform 1 0 2392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 1649977179
transform 1 0 3128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1649977179
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_62
timestamp 1649977179
transform 1 0 6808 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_101
timestamp 1649977179
transform 1 0 10396 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1649977179
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_134
timestamp 1649977179
transform 1 0 13432 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_147
timestamp 1649977179
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1649977179
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_172
timestamp 1649977179
transform 1 0 16928 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_183
timestamp 1649977179
transform 1 0 17940 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1649977179
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_234
timestamp 1649977179
transform 1 0 22632 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_242
timestamp 1649977179
transform 1 0 23368 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_247
timestamp 1649977179
transform 1 0 23828 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1649977179
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_303
timestamp 1649977179
transform 1 0 28980 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_327
timestamp 1649977179
transform 1 0 31188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_357
timestamp 1649977179
transform 1 0 33948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_364
timestamp 1649977179
transform 1 0 34592 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1649977179
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_397
timestamp 1649977179
transform 1 0 37628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_421
timestamp 1649977179
transform 1 0 39836 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_438
timestamp 1649977179
transform 1 0 41400 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1649977179
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_452
timestamp 1649977179
transform 1 0 42688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_459
timestamp 1649977179
transform 1 0 43332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_477
timestamp 1649977179
transform 1 0 44988 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_495
timestamp 1649977179
transform 1 0 46644 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_513
timestamp 1649977179
transform 1 0 48300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_537
timestamp 1649977179
transform 1 0 50508 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_552
timestamp 1649977179
transform 1 0 51888 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_568
timestamp 1649977179
transform 1 0 53360 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_578
timestamp 1649977179
transform 1 0 54280 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_590
timestamp 1649977179
transform 1 0 55384 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_602
timestamp 1649977179
transform 1 0 56488 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_614
timestamp 1649977179
transform 1 0 57592 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1649977179
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_32
timestamp 1649977179
transform 1 0 4048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_56
timestamp 1649977179
transform 1 0 6256 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1649977179
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1649977179
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_110
timestamp 1649977179
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1649977179
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_144
timestamp 1649977179
transform 1 0 14352 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_154
timestamp 1649977179
transform 1 0 15272 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1649977179
transform 1 0 17480 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_201
timestamp 1649977179
transform 1 0 19596 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_212
timestamp 1649977179
transform 1 0 20608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1649977179
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_227
timestamp 1649977179
transform 1 0 21988 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1649977179
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_237
timestamp 1649977179
transform 1 0 22908 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_243
timestamp 1649977179
transform 1 0 23460 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1649977179
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_261
timestamp 1649977179
transform 1 0 25116 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_269
timestamp 1649977179
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_283
timestamp 1649977179
transform 1 0 27140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_290
timestamp 1649977179
transform 1 0 27784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_329
timestamp 1649977179
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_353
timestamp 1649977179
transform 1 0 33580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1649977179
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_378
timestamp 1649977179
transform 1 0 35880 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_386
timestamp 1649977179
transform 1 0 36616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_394
timestamp 1649977179
transform 1 0 37352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_402
timestamp 1649977179
transform 1 0 38088 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_410
timestamp 1649977179
transform 1 0 38824 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_416
timestamp 1649977179
transform 1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_434
timestamp 1649977179
transform 1 0 41032 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_442
timestamp 1649977179
transform 1 0 41768 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_465
timestamp 1649977179
transform 1 0 43884 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_472
timestamp 1649977179
transform 1 0 44528 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_491
timestamp 1649977179
transform 1 0 46276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_497
timestamp 1649977179
transform 1 0 46828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_508
timestamp 1649977179
transform 1 0 47840 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_518
timestamp 1649977179
transform 1 0 48760 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_527
timestamp 1649977179
transform 1 0 49588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_539
timestamp 1649977179
transform 1 0 50692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_546
timestamp 1649977179
transform 1 0 51336 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_571
timestamp 1649977179
transform 1 0 53636 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_579
timestamp 1649977179
transform 1 0 54372 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_596
timestamp 1649977179
transform 1 0 55936 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_602
timestamp 1649977179
transform 1 0 56488 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_607
timestamp 1649977179
transform 1 0 56948 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_619
timestamp 1649977179
transform 1 0 58052 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1649977179
transform 1 0 1748 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_28
timestamp 1649977179
transform 1 0 3680 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1649977179
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_77
timestamp 1649977179
transform 1 0 8188 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_102
timestamp 1649977179
transform 1 0 10488 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1649977179
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_118
timestamp 1649977179
transform 1 0 11960 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_142
timestamp 1649977179
transform 1 0 14168 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_151
timestamp 1649977179
transform 1 0 14996 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_162
timestamp 1649977179
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_179
timestamp 1649977179
transform 1 0 17572 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_187
timestamp 1649977179
transform 1 0 18308 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_192
timestamp 1649977179
transform 1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_196
timestamp 1649977179
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1649977179
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1649977179
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_233
timestamp 1649977179
transform 1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1649977179
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_288
timestamp 1649977179
transform 1 0 27600 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1649977179
transform 1 0 28244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_319
timestamp 1649977179
transform 1 0 30452 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_328
timestamp 1649977179
transform 1 0 31280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1649977179
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_346
timestamp 1649977179
transform 1 0 32936 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_353
timestamp 1649977179
transform 1 0 33580 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_363
timestamp 1649977179
transform 1 0 34500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_377
timestamp 1649977179
transform 1 0 35788 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_396
timestamp 1649977179
transform 1 0 37536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_400
timestamp 1649977179
transform 1 0 37904 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_421
timestamp 1649977179
transform 1 0 39836 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_428
timestamp 1649977179
transform 1 0 40480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_439
timestamp 1649977179
transform 1 0 41492 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_470
timestamp 1649977179
transform 1 0 44344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_495
timestamp 1649977179
transform 1 0 46644 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_510
timestamp 1649977179
transform 1 0 48024 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_534
timestamp 1649977179
transform 1 0 50232 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_548
timestamp 1649977179
transform 1 0 51520 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_565
timestamp 1649977179
transform 1 0 53084 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_577
timestamp 1649977179
transform 1 0 54188 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_589
timestamp 1649977179
transform 1 0 55292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_610
timestamp 1649977179
transform 1 0 57224 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_14
timestamp 1649977179
transform 1 0 2392 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_20
timestamp 1649977179
transform 1 0 2944 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_32
timestamp 1649977179
transform 1 0 4048 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_56
timestamp 1649977179
transform 1 0 6256 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1649977179
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1649977179
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1649977179
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1649977179
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_161
timestamp 1649977179
transform 1 0 15916 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_168
timestamp 1649977179
transform 1 0 16560 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1649977179
transform 1 0 17572 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_204
timestamp 1649977179
transform 1 0 19872 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_208
timestamp 1649977179
transform 1 0 20240 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1649977179
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_219
timestamp 1649977179
transform 1 0 21252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_228
timestamp 1649977179
transform 1 0 22080 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_238
timestamp 1649977179
transform 1 0 23000 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_259
timestamp 1649977179
transform 1 0 24932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_263
timestamp 1649977179
transform 1 0 25300 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_267
timestamp 1649977179
transform 1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_275
timestamp 1649977179
transform 1 0 26404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_279
timestamp 1649977179
transform 1 0 26772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_283
timestamp 1649977179
transform 1 0 27140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_295
timestamp 1649977179
transform 1 0 28244 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1649977179
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_315
timestamp 1649977179
transform 1 0 30084 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_322
timestamp 1649977179
transform 1 0 30728 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_326
timestamp 1649977179
transform 1 0 31096 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_340
timestamp 1649977179
transform 1 0 32384 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_352
timestamp 1649977179
transform 1 0 33488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_356
timestamp 1649977179
transform 1 0 33856 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1649977179
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_369
timestamp 1649977179
transform 1 0 35052 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_383
timestamp 1649977179
transform 1 0 36340 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_407
timestamp 1649977179
transform 1 0 38548 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_415
timestamp 1649977179
transform 1 0 39284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_424
timestamp 1649977179
transform 1 0 40112 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_436
timestamp 1649977179
transform 1 0 41216 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_448
timestamp 1649977179
transform 1 0 42320 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_460
timestamp 1649977179
transform 1 0 43424 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_465
timestamp 1649977179
transform 1 0 43884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1649977179
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_484
timestamp 1649977179
transform 1 0 45632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_490
timestamp 1649977179
transform 1 0 46184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_496
timestamp 1649977179
transform 1 0 46736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_502
timestamp 1649977179
transform 1 0 47288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_506
timestamp 1649977179
transform 1 0 47656 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_517
timestamp 1649977179
transform 1 0 48668 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_528
timestamp 1649977179
transform 1 0 49680 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_535
timestamp 1649977179
transform 1 0 50324 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_546
timestamp 1649977179
transform 1 0 51336 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_570
timestamp 1649977179
transform 1 0 53544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_582
timestamp 1649977179
transform 1 0 54648 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_593
timestamp 1649977179
transform 1 0 55660 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_605
timestamp 1649977179
transform 1 0 56764 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_617
timestamp 1649977179
transform 1 0 57868 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_7
timestamp 1649977179
transform 1 0 1748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_30
timestamp 1649977179
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_34
timestamp 1649977179
transform 1 0 4232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_38
timestamp 1649977179
transform 1 0 4600 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_45
timestamp 1649977179
transform 1 0 5244 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1649977179
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_84
timestamp 1649977179
transform 1 0 8832 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1649977179
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_117
timestamp 1649977179
transform 1 0 11868 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1649977179
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_133
timestamp 1649977179
transform 1 0 13340 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_157
timestamp 1649977179
transform 1 0 15548 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1649977179
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_173
timestamp 1649977179
transform 1 0 17020 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1649977179
transform 1 0 17572 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_213
timestamp 1649977179
transform 1 0 20700 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1649977179
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1649977179
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_242
timestamp 1649977179
transform 1 0 23368 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_246
timestamp 1649977179
transform 1 0 23736 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_253
timestamp 1649977179
transform 1 0 24380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_264
timestamp 1649977179
transform 1 0 25392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 1649977179
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_289
timestamp 1649977179
transform 1 0 27692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_303
timestamp 1649977179
transform 1 0 28980 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_311
timestamp 1649977179
transform 1 0 29716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1649977179
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_340
timestamp 1649977179
transform 1 0 32384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_344
timestamp 1649977179
transform 1 0 32752 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_348
timestamp 1649977179
transform 1 0 33120 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_356
timestamp 1649977179
transform 1 0 33856 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_378
timestamp 1649977179
transform 1 0 35880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_397
timestamp 1649977179
transform 1 0 37628 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_401
timestamp 1649977179
transform 1 0 37996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_408
timestamp 1649977179
transform 1 0 38640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_412
timestamp 1649977179
transform 1 0 39008 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_416
timestamp 1649977179
transform 1 0 39376 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_428
timestamp 1649977179
transform 1 0 40480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1649977179
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_451
timestamp 1649977179
transform 1 0 42596 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_463
timestamp 1649977179
transform 1 0 43700 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_476
timestamp 1649977179
transform 1 0 44896 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1649977179
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_507
timestamp 1649977179
transform 1 0 47748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_532
timestamp 1649977179
transform 1 0 50048 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_540
timestamp 1649977179
transform 1 0 50784 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_548
timestamp 1649977179
transform 1 0 51520 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_554
timestamp 1649977179
transform 1 0 52072 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_6
timestamp 1649977179
transform 1 0 1656 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_13
timestamp 1649977179
transform 1 0 2300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1649977179
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_50
timestamp 1649977179
transform 1 0 5704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_58
timestamp 1649977179
transform 1 0 6440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1649977179
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_88
timestamp 1649977179
transform 1 0 9200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_112
timestamp 1649977179
transform 1 0 11408 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1649977179
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_161
timestamp 1649977179
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_169
timestamp 1649977179
transform 1 0 16652 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_180
timestamp 1649977179
transform 1 0 17664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_205
timestamp 1649977179
transform 1 0 19964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_211
timestamp 1649977179
transform 1 0 20516 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_230
timestamp 1649977179
transform 1 0 22264 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_238
timestamp 1649977179
transform 1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_242
timestamp 1649977179
transform 1 0 23368 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1649977179
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_261
timestamp 1649977179
transform 1 0 25116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_272
timestamp 1649977179
transform 1 0 26128 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_282
timestamp 1649977179
transform 1 0 27048 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 1649977179
transform 1 0 27600 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1649977179
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_319
timestamp 1649977179
transform 1 0 30452 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_325
timestamp 1649977179
transform 1 0 31004 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_346
timestamp 1649977179
transform 1 0 32936 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_354
timestamp 1649977179
transform 1 0 33672 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1649977179
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_374
timestamp 1649977179
transform 1 0 35512 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_381
timestamp 1649977179
transform 1 0 36156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_393
timestamp 1649977179
transform 1 0 37260 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_405
timestamp 1649977179
transform 1 0 38364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_417
timestamp 1649977179
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_460
timestamp 1649977179
transform 1 0 43424 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1649977179
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_491
timestamp 1649977179
transform 1 0 46276 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_497
timestamp 1649977179
transform 1 0 46828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_503
timestamp 1649977179
transform 1 0 47380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_528
timestamp 1649977179
transform 1 0 49680 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_6
timestamp 1649977179
transform 1 0 1656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1649977179
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_25
timestamp 1649977179
transform 1 0 3404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_36
timestamp 1649977179
transform 1 0 4416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_43
timestamp 1649977179
transform 1 0 5060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1649977179
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_60
timestamp 1649977179
transform 1 0 6624 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_84
timestamp 1649977179
transform 1 0 8832 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1649977179
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1649977179
transform 1 0 13524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_159
timestamp 1649977179
transform 1 0 15732 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_173
timestamp 1649977179
transform 1 0 17020 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_186
timestamp 1649977179
transform 1 0 18216 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_194
timestamp 1649977179
transform 1 0 18952 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_198
timestamp 1649977179
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_212
timestamp 1649977179
transform 1 0 20608 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_216
timestamp 1649977179
transform 1 0 20976 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1649977179
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_235
timestamp 1649977179
transform 1 0 22724 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_251
timestamp 1649977179
transform 1 0 24196 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_260
timestamp 1649977179
transform 1 0 25024 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1649977179
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_285
timestamp 1649977179
transform 1 0 27324 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_302
timestamp 1649977179
transform 1 0 28888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_313
timestamp 1649977179
transform 1 0 29900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_321
timestamp 1649977179
transform 1 0 30636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_328
timestamp 1649977179
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_340
timestamp 1649977179
transform 1 0 32384 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_352
timestamp 1649977179
transform 1 0 33488 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_374
timestamp 1649977179
transform 1 0 35512 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_386
timestamp 1649977179
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_413
timestamp 1649977179
transform 1 0 39100 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_430
timestamp 1649977179
transform 1 0 40664 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_442
timestamp 1649977179
transform 1 0 41768 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_526
timestamp 1649977179
transform 1 0 49496 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_538
timestamp 1649977179
transform 1 0 50600 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_550
timestamp 1649977179
transform 1 0 51704 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_558
timestamp 1649977179
transform 1 0 52440 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_621
timestamp 1649977179
transform 1 0 58236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1649977179
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_32
timestamp 1649977179
transform 1 0 4048 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_36
timestamp 1649977179
transform 1 0 4416 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_67
timestamp 1649977179
transform 1 0 7268 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1649977179
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_89
timestamp 1649977179
transform 1 0 9292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp 1649977179
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_150
timestamp 1649977179
transform 1 0 14904 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_158
timestamp 1649977179
transform 1 0 15640 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1649977179
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_227
timestamp 1649977179
transform 1 0 21988 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_237
timestamp 1649977179
transform 1 0 22908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1649977179
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_255
timestamp 1649977179
transform 1 0 24564 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_261
timestamp 1649977179
transform 1 0 25116 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_272
timestamp 1649977179
transform 1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_296
timestamp 1649977179
transform 1 0 28336 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_300
timestamp 1649977179
transform 1 0 28704 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1649977179
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_339
timestamp 1649977179
transform 1 0 32292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1649977179
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_380
timestamp 1649977179
transform 1 0 36064 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_387
timestamp 1649977179
transform 1 0 36708 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_399
timestamp 1649977179
transform 1 0 37812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_403
timestamp 1649977179
transform 1 0 38180 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_407
timestamp 1649977179
transform 1 0 38548 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_414
timestamp 1649977179
transform 1 0 39192 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_424
timestamp 1649977179
transform 1 0 40112 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_436
timestamp 1649977179
transform 1 0 41216 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_448
timestamp 1649977179
transform 1 0 42320 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_460
timestamp 1649977179
transform 1 0 43424 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_472
timestamp 1649977179
transform 1 0 44528 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_507
timestamp 1649977179
transform 1 0 47748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_519
timestamp 1649977179
transform 1 0 48852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_7
timestamp 1649977179
transform 1 0 1748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_10
timestamp 1649977179
transform 1 0 2024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_16
timestamp 1649977179
transform 1 0 2576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_22
timestamp 1649977179
transform 1 0 3128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_33
timestamp 1649977179
transform 1 0 4140 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_37
timestamp 1649977179
transform 1 0 4508 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_41
timestamp 1649977179
transform 1 0 4876 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1649977179
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_126
timestamp 1649977179
transform 1 0 12696 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_136
timestamp 1649977179
transform 1 0 13616 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_143
timestamp 1649977179
transform 1 0 14260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_154
timestamp 1649977179
transform 1 0 15272 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_160
timestamp 1649977179
transform 1 0 15824 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1649977179
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_173
timestamp 1649977179
transform 1 0 17020 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_187
timestamp 1649977179
transform 1 0 18308 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_194
timestamp 1649977179
transform 1 0 18952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1649977179
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_228
timestamp 1649977179
transform 1 0 22080 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_242
timestamp 1649977179
transform 1 0 23368 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_253
timestamp 1649977179
transform 1 0 24380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_267
timestamp 1649977179
transform 1 0 25668 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1649977179
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_287
timestamp 1649977179
transform 1 0 27508 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_298
timestamp 1649977179
transform 1 0 28520 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_302
timestamp 1649977179
transform 1 0 28888 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_306
timestamp 1649977179
transform 1 0 29256 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_310
timestamp 1649977179
transform 1 0 29624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_315
timestamp 1649977179
transform 1 0 30084 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1649977179
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_380
timestamp 1649977179
transform 1 0 36064 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_414
timestamp 1649977179
transform 1 0 39192 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_426
timestamp 1649977179
transform 1 0 40296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_438
timestamp 1649977179
transform 1 0 41400 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1649977179
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_7
timestamp 1649977179
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_11
timestamp 1649977179
transform 1 0 2116 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_21
timestamp 1649977179
transform 1 0 3036 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1649977179
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_50
timestamp 1649977179
transform 1 0 5704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_56
timestamp 1649977179
transform 1 0 6256 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_67
timestamp 1649977179
transform 1 0 7268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1649977179
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_89
timestamp 1649977179
transform 1 0 9292 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_93
timestamp 1649977179
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1649977179
transform 1 0 10396 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_112
timestamp 1649977179
transform 1 0 11408 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_118
timestamp 1649977179
transform 1 0 11960 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_126
timestamp 1649977179
transform 1 0 12696 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_151
timestamp 1649977179
transform 1 0 14996 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_159
timestamp 1649977179
transform 1 0 15732 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_163
timestamp 1649977179
transform 1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_174
timestamp 1649977179
transform 1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_185
timestamp 1649977179
transform 1 0 18124 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1649977179
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_204
timestamp 1649977179
transform 1 0 19872 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_230
timestamp 1649977179
transform 1 0 22264 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_236
timestamp 1649977179
transform 1 0 22816 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_239
timestamp 1649977179
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_273
timestamp 1649977179
transform 1 0 26220 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_294
timestamp 1649977179
transform 1 0 28152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_329
timestamp 1649977179
transform 1 0 31372 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_336
timestamp 1649977179
transform 1 0 32016 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_348
timestamp 1649977179
transform 1 0 33120 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1649977179
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_369
timestamp 1649977179
transform 1 0 35052 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_381
timestamp 1649977179
transform 1 0 36156 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_393
timestamp 1649977179
transform 1 0 37260 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_405
timestamp 1649977179
transform 1 0 38364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_417
timestamp 1649977179
transform 1 0 39468 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_23
timestamp 1649977179
transform 1 0 3220 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_32
timestamp 1649977179
transform 1 0 4048 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_38
timestamp 1649977179
transform 1 0 4600 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_46
timestamp 1649977179
transform 1 0 5336 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1649977179
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_68
timestamp 1649977179
transform 1 0 7360 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_77
timestamp 1649977179
transform 1 0 8188 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_84
timestamp 1649977179
transform 1 0 8832 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1649977179
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_120
timestamp 1649977179
transform 1 0 12144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_126
timestamp 1649977179
transform 1 0 12696 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_134
timestamp 1649977179
transform 1 0 13432 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1649977179
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1649977179
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_179
timestamp 1649977179
transform 1 0 17572 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_183
timestamp 1649977179
transform 1 0 17940 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_204
timestamp 1649977179
transform 1 0 19872 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_215
timestamp 1649977179
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_232
timestamp 1649977179
transform 1 0 22448 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_248
timestamp 1649977179
transform 1 0 23920 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_260
timestamp 1649977179
transform 1 0 25024 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_272
timestamp 1649977179
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1649977179
transform 1 0 28244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_319
timestamp 1649977179
transform 1 0 30452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_326
timestamp 1649977179
transform 1 0 31096 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1649977179
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_11
timestamp 1649977179
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_21
timestamp 1649977179
transform 1 0 3036 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1649977179
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_49
timestamp 1649977179
transform 1 0 5612 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_62
timestamp 1649977179
transform 1 0 6808 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1649977179
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_89
timestamp 1649977179
transform 1 0 9292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_129
timestamp 1649977179
transform 1 0 12972 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1649977179
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1649977179
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_161
timestamp 1649977179
transform 1 0 15916 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_167
timestamp 1649977179
transform 1 0 16468 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_172
timestamp 1649977179
transform 1 0 16928 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_181
timestamp 1649977179
transform 1 0 17756 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_187
timestamp 1649977179
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1649977179
transform 1 0 20056 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_214
timestamp 1649977179
transform 1 0 20792 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_226
timestamp 1649977179
transform 1 0 21896 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1649977179
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_261
timestamp 1649977179
transform 1 0 25116 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_273
timestamp 1649977179
transform 1 0 26220 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_285
timestamp 1649977179
transform 1 0 27324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1649977179
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1649977179
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_406
timestamp 1649977179
transform 1 0 38456 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_418
timestamp 1649977179
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_17
timestamp 1649977179
transform 1 0 2668 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_25
timestamp 1649977179
transform 1 0 3404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_32
timestamp 1649977179
transform 1 0 4048 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_40
timestamp 1649977179
transform 1 0 4784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 1649977179
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1649977179
transform 1 0 8188 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1649977179
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_90
timestamp 1649977179
transform 1 0 9384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_102
timestamp 1649977179
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1649977179
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_115
timestamp 1649977179
transform 1 0 11684 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_123
timestamp 1649977179
transform 1 0 12420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_148
timestamp 1649977179
transform 1 0 14720 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_156
timestamp 1649977179
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_172
timestamp 1649977179
transform 1 0 16928 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_178
timestamp 1649977179
transform 1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_185
timestamp 1649977179
transform 1 0 18124 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_200
timestamp 1649977179
transform 1 0 19504 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_206
timestamp 1649977179
transform 1 0 20056 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_218
timestamp 1649977179
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_241
timestamp 1649977179
transform 1 0 23276 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_246
timestamp 1649977179
transform 1 0 23736 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_252
timestamp 1649977179
transform 1 0 24288 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_264
timestamp 1649977179
transform 1 0 25392 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1649977179
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1649977179
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_35
timestamp 1649977179
transform 1 0 4324 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_43
timestamp 1649977179
transform 1 0 5060 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_47
timestamp 1649977179
transform 1 0 5428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_59
timestamp 1649977179
transform 1 0 6532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_71
timestamp 1649977179
transform 1 0 7636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_79
timestamp 1649977179
transform 1 0 8372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_98
timestamp 1649977179
transform 1 0 10120 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_110
timestamp 1649977179
transform 1 0 11224 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_122
timestamp 1649977179
transform 1 0 12328 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 1649977179
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_155
timestamp 1649977179
transform 1 0 15364 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_179
timestamp 1649977179
transform 1 0 17572 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1649977179
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_210
timestamp 1649977179
transform 1 0 20424 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_222
timestamp 1649977179
transform 1 0 21528 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_234
timestamp 1649977179
transform 1 0 22632 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_246
timestamp 1649977179
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_370
timestamp 1649977179
transform 1 0 35144 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_382
timestamp 1649977179
transform 1 0 36248 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_394
timestamp 1649977179
transform 1 0 37352 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_406
timestamp 1649977179
transform 1 0 38456 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1649977179
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_621
timestamp 1649977179
transform 1 0 58236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_9
timestamp 1649977179
transform 1 0 1932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_33
timestamp 1649977179
transform 1 0 4140 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1649977179
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_64
timestamp 1649977179
transform 1 0 6992 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_72
timestamp 1649977179
transform 1 0 7728 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_79
timestamp 1649977179
transform 1 0 8372 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_98
timestamp 1649977179
transform 1 0 10120 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1649977179
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_173
timestamp 1649977179
transform 1 0 17020 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_179
timestamp 1649977179
transform 1 0 17572 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_187
timestamp 1649977179
transform 1 0 18308 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_213
timestamp 1649977179
transform 1 0 20700 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1649977179
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_366
timestamp 1649977179
transform 1 0 34776 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1649977179
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_621
timestamp 1649977179
transform 1 0 58236 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_39
timestamp 1649977179
transform 1 0 4692 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_49
timestamp 1649977179
transform 1 0 5612 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_60
timestamp 1649977179
transform 1 0 6624 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_78
timestamp 1649977179
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_87
timestamp 1649977179
transform 1 0 9108 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_93
timestamp 1649977179
transform 1 0 9660 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_105
timestamp 1649977179
transform 1 0 10764 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_117
timestamp 1649977179
transform 1 0 11868 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_129
timestamp 1649977179
transform 1 0 12972 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1649977179
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_149
timestamp 1649977179
transform 1 0 14812 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_161
timestamp 1649977179
transform 1 0 15916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_173
timestamp 1649977179
transform 1 0 17020 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_181
timestamp 1649977179
transform 1 0 17756 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_186
timestamp 1649977179
transform 1 0 18216 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1649977179
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_201
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_213
timestamp 1649977179
transform 1 0 20700 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_225
timestamp 1649977179
transform 1 0 21804 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_237
timestamp 1649977179
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1649977179
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_281
timestamp 1649977179
transform 1 0 26956 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_288
timestamp 1649977179
transform 1 0 27600 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_300
timestamp 1649977179
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1649977179
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_383
timestamp 1649977179
transform 1 0 36340 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_395
timestamp 1649977179
transform 1 0 37444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_407
timestamp 1649977179
transform 1 0 38548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_11
timestamp 1649977179
transform 1 0 2116 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_35
timestamp 1649977179
transform 1 0 4324 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_41
timestamp 1649977179
transform 1 0 4876 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_48
timestamp 1649977179
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_77
timestamp 1649977179
transform 1 0 8188 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_85
timestamp 1649977179
transform 1 0 8924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_97
timestamp 1649977179
transform 1 0 10028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1649977179
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_177
timestamp 1649977179
transform 1 0 17388 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_195
timestamp 1649977179
transform 1 0 19044 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_201
timestamp 1649977179
transform 1 0 19596 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_215
timestamp 1649977179
transform 1 0 20884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_252
timestamp 1649977179
transform 1 0 24288 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1649977179
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_295
timestamp 1649977179
transform 1 0 28244 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_307
timestamp 1649977179
transform 1 0 29348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_319
timestamp 1649977179
transform 1 0 30452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1649977179
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_367
timestamp 1649977179
transform 1 0 34868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_379
timestamp 1649977179
transform 1 0 35972 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1649977179
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_21
timestamp 1649977179
transform 1 0 3036 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1649977179
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_49
timestamp 1649977179
transform 1 0 5612 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_56
timestamp 1649977179
transform 1 0 6256 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_68
timestamp 1649977179
transform 1 0 7360 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_76
timestamp 1649977179
transform 1 0 8096 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_79
timestamp 1649977179
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_152
timestamp 1649977179
transform 1 0 15088 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_160
timestamp 1649977179
transform 1 0 15824 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_184
timestamp 1649977179
transform 1 0 18032 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_217
timestamp 1649977179
transform 1 0 21068 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_229
timestamp 1649977179
transform 1 0 22172 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1649977179
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1649977179
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_273
timestamp 1649977179
transform 1 0 26220 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_276
timestamp 1649977179
transform 1 0 26496 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1649977179
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_311
timestamp 1649977179
transform 1 0 29716 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_323
timestamp 1649977179
transform 1 0 30820 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_335
timestamp 1649977179
transform 1 0 31924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_347
timestamp 1649977179
transform 1 0 33028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1649977179
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_373
timestamp 1649977179
transform 1 0 35420 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_376
timestamp 1649977179
transform 1 0 35696 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_394
timestamp 1649977179
transform 1 0 37352 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_406
timestamp 1649977179
transform 1 0 38456 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_418
timestamp 1649977179
transform 1 0 39560 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_31
timestamp 1649977179
transform 1 0 3956 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_34
timestamp 1649977179
transform 1 0 4232 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1649977179
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_60
timestamp 1649977179
transform 1 0 6624 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_66
timestamp 1649977179
transform 1 0 7176 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_72
timestamp 1649977179
transform 1 0 7728 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_78
timestamp 1649977179
transform 1 0 8280 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_90
timestamp 1649977179
transform 1 0 9384 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_102
timestamp 1649977179
transform 1 0 10488 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1649977179
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_145
timestamp 1649977179
transform 1 0 14444 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_155
timestamp 1649977179
transform 1 0 15364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_197
timestamp 1649977179
transform 1 0 19228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_202
timestamp 1649977179
transform 1 0 19688 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_214
timestamp 1649977179
transform 1 0 20792 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1649977179
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_377
timestamp 1649977179
transform 1 0 35788 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_380
timestamp 1649977179
transform 1 0 36064 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_396
timestamp 1649977179
transform 1 0 37536 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_402
timestamp 1649977179
transform 1 0 38088 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_414
timestamp 1649977179
transform 1 0 39192 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_426
timestamp 1649977179
transform 1 0 40296 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_438
timestamp 1649977179
transform 1 0 41400 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_446
timestamp 1649977179
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_7
timestamp 1649977179
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_11
timestamp 1649977179
transform 1 0 2116 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1649977179
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_37
timestamp 1649977179
transform 1 0 4508 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_40
timestamp 1649977179
transform 1 0 4784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_58
timestamp 1649977179
transform 1 0 6440 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_76
timestamp 1649977179
transform 1 0 8096 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_87
timestamp 1649977179
transform 1 0 9108 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_99
timestamp 1649977179
transform 1 0 10212 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_111
timestamp 1649977179
transform 1 0 11316 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_123
timestamp 1649977179
transform 1 0 12420 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_135
timestamp 1649977179
transform 1 0 13524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_370
timestamp 1649977179
transform 1 0 35144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_376
timestamp 1649977179
transform 1 0 35696 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_394
timestamp 1649977179
transform 1 0 37352 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_412
timestamp 1649977179
transform 1 0 39008 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_31
timestamp 1649977179
transform 1 0 3956 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_34
timestamp 1649977179
transform 1 0 4232 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1649977179
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_71
timestamp 1649977179
transform 1 0 7636 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_77
timestamp 1649977179
transform 1 0 8188 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_83
timestamp 1649977179
transform 1 0 8740 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_95
timestamp 1649977179
transform 1 0 9844 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1649977179
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_367
timestamp 1649977179
transform 1 0 34868 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_370
timestamp 1649977179
transform 1 0 35144 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1649977179
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_407
timestamp 1649977179
transform 1 0 38548 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_413
timestamp 1649977179
transform 1 0 39100 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_419
timestamp 1649977179
transform 1 0 39652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_431
timestamp 1649977179
transform 1 0 40756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_443
timestamp 1649977179
transform 1 0 41860 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_489
timestamp 1649977179
transform 1 0 46092 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_495
timestamp 1649977179
transform 1 0 46644 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_23
timestamp 1649977179
transform 1 0 3220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_37
timestamp 1649977179
transform 1 0 4508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_40
timestamp 1649977179
transform 1 0 4784 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_58
timestamp 1649977179
transform 1 0 6440 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_76
timestamp 1649977179
transform 1 0 8096 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_87
timestamp 1649977179
transform 1 0 9108 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_93
timestamp 1649977179
transform 1 0 9660 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_105
timestamp 1649977179
transform 1 0 10764 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_117
timestamp 1649977179
transform 1 0 11868 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_129
timestamp 1649977179
transform 1 0 12972 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_137
timestamp 1649977179
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_371
timestamp 1649977179
transform 1 0 35236 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_374
timestamp 1649977179
transform 1 0 35512 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_394
timestamp 1649977179
transform 1 0 37352 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_412
timestamp 1649977179
transform 1 0 39008 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_21
timestamp 1649977179
transform 1 0 3036 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_35
timestamp 1649977179
transform 1 0 4324 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_40
timestamp 1649977179
transform 1 0 4784 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_48
timestamp 1649977179
transform 1 0 5520 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1649977179
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_60
timestamp 1649977179
transform 1 0 6624 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_87
timestamp 1649977179
transform 1 0 9108 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_378
timestamp 1649977179
transform 1 0 35880 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_384
timestamp 1649977179
transform 1 0 36432 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_396
timestamp 1649977179
transform 1 0 37536 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1649977179
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_409
timestamp 1649977179
transform 1 0 38732 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_415
timestamp 1649977179
transform 1 0 39284 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_427
timestamp 1649977179
transform 1 0 40388 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_439
timestamp 1649977179
transform 1 0 41492 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_38
timestamp 1649977179
transform 1 0 4600 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_58
timestamp 1649977179
transform 1 0 6440 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_64
timestamp 1649977179
transform 1 0 6992 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_70
timestamp 1649977179
transform 1 0 7544 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1649977179
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1649977179
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_201
timestamp 1649977179
transform 1 0 19596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_213
timestamp 1649977179
transform 1 0 20700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_225
timestamp 1649977179
transform 1 0 21804 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_238
timestamp 1649977179
transform 1 0 23000 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_244
timestamp 1649977179
transform 1 0 23552 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_342
timestamp 1649977179
transform 1 0 32568 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_348
timestamp 1649977179
transform 1 0 33120 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1649977179
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_373
timestamp 1649977179
transform 1 0 35420 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_376
timestamp 1649977179
transform 1 0 35696 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_394
timestamp 1649977179
transform 1 0 37352 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_402
timestamp 1649977179
transform 1 0 38088 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_414
timestamp 1649977179
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_424
timestamp 1649977179
transform 1 0 40112 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_436
timestamp 1649977179
transform 1 0 41216 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_448
timestamp 1649977179
transform 1 0 42320 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_460
timestamp 1649977179
transform 1 0 43424 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_472
timestamp 1649977179
transform 1 0 44528 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_563
timestamp 1649977179
transform 1 0 52900 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_575
timestamp 1649977179
transform 1 0 54004 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_609
timestamp 1649977179
transform 1 0 57132 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_614
timestamp 1649977179
transform 1 0 57592 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_622
timestamp 1649977179
transform 1 0 58328 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_7
timestamp 1649977179
transform 1 0 1748 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_19
timestamp 1649977179
transform 1 0 2852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_29
timestamp 1649977179
transform 1 0 3772 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_37
timestamp 1649977179
transform 1 0 4508 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_42
timestamp 1649977179
transform 1 0 4968 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1649977179
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_62
timestamp 1649977179
transform 1 0 6808 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_68
timestamp 1649977179
transform 1 0 7360 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_80
timestamp 1649977179
transform 1 0 8464 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_85
timestamp 1649977179
transform 1 0 8924 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_91
timestamp 1649977179
transform 1 0 9476 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_103
timestamp 1649977179
transform 1 0 10580 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_141
timestamp 1649977179
transform 1 0 14076 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_147
timestamp 1649977179
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_159
timestamp 1649977179
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_200
timestamp 1649977179
transform 1 0 19504 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_212
timestamp 1649977179
transform 1 0 20608 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_256
timestamp 1649977179
transform 1 0 24656 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_262
timestamp 1649977179
transform 1 0 25208 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_274
timestamp 1649977179
transform 1 0 26312 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_289
timestamp 1649977179
transform 1 0 27692 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_301
timestamp 1649977179
transform 1 0 28796 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_307
timestamp 1649977179
transform 1 0 29348 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_309
timestamp 1649977179
transform 1 0 29532 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_357
timestamp 1649977179
transform 1 0 33948 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_363
timestamp 1649977179
transform 1 0 34500 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_365
timestamp 1649977179
transform 1 0 34684 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_377
timestamp 1649977179
transform 1 0 35788 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_380
timestamp 1649977179
transform 1 0 36064 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_398
timestamp 1649977179
transform 1 0 37720 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_406
timestamp 1649977179
transform 1 0 38456 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_412
timestamp 1649977179
transform 1 0 39008 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_421
timestamp 1649977179
transform 1 0 39836 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_433
timestamp 1649977179
transform 1 0 40940 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_445
timestamp 1649977179
transform 1 0 42044 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_457
timestamp 1649977179
transform 1 0 43148 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_477
timestamp 1649977179
transform 1 0 44988 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_489
timestamp 1649977179
transform 1 0 46092 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_501
timestamp 1649977179
transform 1 0 47196 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_513
timestamp 1649977179
transform 1 0 48300 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_518
timestamp 1649977179
transform 1 0 48760 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_530
timestamp 1649977179
transform 1 0 49864 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_533
timestamp 1649977179
transform 1 0 50140 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_545
timestamp 1649977179
transform 1 0 51244 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_557
timestamp 1649977179
transform 1 0 52348 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_567
timestamp 1649977179
transform 1 0 53268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_579
timestamp 1649977179
transform 1 0 54372 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_587
timestamp 1649977179
transform 1 0 55108 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_589
timestamp 1649977179
transform 1 0 55292 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_601
timestamp 1649977179
transform 1 0 56396 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_612
timestamp 1649977179
transform 1 0 57408 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1649977179
transform 1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 3680 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 8832 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 13984 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 19136 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 24288 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 29440 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 34592 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 39744 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 44896 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 50048 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 55200 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0485__1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 34224 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0486_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23000 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0487_
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0488__6
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0489__7
timestamp 1649977179
transform -1 0 24656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0490__8
timestamp 1649977179
transform -1 0 24932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491__9
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492__10
timestamp 1649977179
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0493_
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494__11
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0495__12
timestamp 1649977179
transform -1 0 25668 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0496__13
timestamp 1649977179
transform -1 0 23920 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0497__14
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0498__15
timestamp 1649977179
transform 1 0 22356 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0499_
timestamp 1649977179
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0500_
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0501__16
timestamp 1649977179
transform -1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0502__17
timestamp 1649977179
transform -1 0 14076 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0503__18
timestamp 1649977179
transform -1 0 12604 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0504__19
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0505__20
timestamp 1649977179
transform -1 0 12604 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0506_
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0507__21
timestamp 1649977179
transform 1 0 5612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0508__22
timestamp 1649977179
transform -1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0509__23
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0510__24
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0511_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35788 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0512_
timestamp 1649977179
transform -1 0 34592 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0513_
timestamp 1649977179
transform -1 0 38180 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _0514_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 38088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0515_
timestamp 1649977179
transform 1 0 38916 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0516_
timestamp 1649977179
transform -1 0 28796 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0517_
timestamp 1649977179
transform -1 0 31096 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0518_
timestamp 1649977179
transform -1 0 36064 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0519_
timestamp 1649977179
transform 1 0 37720 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0520_
timestamp 1649977179
transform 1 0 38456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0521_
timestamp 1649977179
transform 1 0 40940 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0522_
timestamp 1649977179
transform -1 0 31004 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0523_
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0524_
timestamp 1649977179
transform 1 0 40848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0526_
timestamp 1649977179
transform -1 0 36616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0527_
timestamp 1649977179
transform -1 0 36156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1649977179
transform -1 0 25668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1649977179
transform -1 0 32384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0532_
timestamp 1649977179
transform -1 0 36340 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1649977179
transform 1 0 38548 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1649977179
transform -1 0 29808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1649977179
transform -1 0 27784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1649977179
transform -1 0 37168 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537__25
timestamp 1649977179
transform 1 0 6532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0538_
timestamp 1649977179
transform -1 0 5244 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0539__26
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0540__27
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0541__28
timestamp 1649977179
transform -1 0 3312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0542_
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0543_
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0544_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10120 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  _0545_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0546_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3496 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0547_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0548_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6992 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0549_
timestamp 1649977179
transform -1 0 6808 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1649977179
transform -1 0 3220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0551_
timestamp 1649977179
transform -1 0 2484 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _0552_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0553_
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0554_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4048 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0555_
timestamp 1649977179
transform -1 0 2392 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0556_
timestamp 1649977179
transform -1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0557_
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0558_
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0559_
timestamp 1649977179
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0560_
timestamp 1649977179
transform 1 0 16928 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0561_
timestamp 1649977179
transform 1 0 22632 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0562_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0563_
timestamp 1649977179
transform -1 0 9292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0564_
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0565_
timestamp 1649977179
transform 1 0 20240 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0566_
timestamp 1649977179
transform -1 0 19320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0567_
timestamp 1649977179
transform -1 0 23644 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0568_
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0569_
timestamp 1649977179
transform -1 0 23920 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0570_
timestamp 1649977179
transform 1 0 19228 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1649977179
transform -1 0 18768 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0572_
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_4  _0573_
timestamp 1649977179
transform 1 0 5244 0 1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__or4b_1  _0574_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18032 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0575_
timestamp 1649977179
transform 1 0 9660 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0576_
timestamp 1649977179
transform 1 0 12604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _0577_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1649977179
transform 1 0 13064 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0579_
timestamp 1649977179
transform 1 0 15272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0580_
timestamp 1649977179
transform 1 0 16560 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _0581_
timestamp 1649977179
transform 1 0 16192 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0582_
timestamp 1649977179
transform 1 0 23736 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0583_
timestamp 1649977179
transform -1 0 23368 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0584_
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0585_
timestamp 1649977179
transform 1 0 20424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0586_
timestamp 1649977179
transform -1 0 18216 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0587_
timestamp 1649977179
transform 1 0 19688 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0588_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20608 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0589_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0590_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17020 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0591_
timestamp 1649977179
transform -1 0 5888 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0592_
timestamp 1649977179
transform -1 0 7360 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0593_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3404 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0594_
timestamp 1649977179
transform -1 0 3312 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0595_
timestamp 1649977179
transform 1 0 3772 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0596_
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0597_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18952 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0598_
timestamp 1649977179
transform -1 0 20608 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0599_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0600_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5428 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0601_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0602_
timestamp 1649977179
transform -1 0 8280 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0603_
timestamp 1649977179
transform 1 0 6624 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0604_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0605_
timestamp 1649977179
transform -1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0606_
timestamp 1649977179
transform 1 0 20976 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0607_
timestamp 1649977179
transform 1 0 17940 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0608_
timestamp 1649977179
transform -1 0 11408 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0609_
timestamp 1649977179
transform -1 0 13248 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0610_
timestamp 1649977179
transform -1 0 29072 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0611_
timestamp 1649977179
transform -1 0 22080 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0612_
timestamp 1649977179
transform -1 0 21344 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0613_
timestamp 1649977179
transform 1 0 19412 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0614_
timestamp 1649977179
transform 1 0 22080 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0615_
timestamp 1649977179
transform -1 0 14720 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0616_
timestamp 1649977179
transform -1 0 14996 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0617_
timestamp 1649977179
transform -1 0 16192 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0618_
timestamp 1649977179
transform 1 0 22448 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0619_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23736 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0620_
timestamp 1649977179
transform 1 0 16468 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0621_
timestamp 1649977179
transform -1 0 17756 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0622_
timestamp 1649977179
transform -1 0 21252 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0623_
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0624_
timestamp 1649977179
transform -1 0 19872 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0625_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17020 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0626_
timestamp 1649977179
transform 1 0 21160 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _0627_
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__clkinv_2  _0628_
timestamp 1649977179
transform 1 0 32384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0629_
timestamp 1649977179
transform -1 0 20608 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0630_
timestamp 1649977179
transform 1 0 18308 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0631_
timestamp 1649977179
transform -1 0 16008 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0632_
timestamp 1649977179
transform -1 0 14996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0633_
timestamp 1649977179
transform -1 0 28336 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0634_
timestamp 1649977179
transform 1 0 20148 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1649977179
transform 1 0 27324 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0636_
timestamp 1649977179
transform 1 0 20240 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0637_
timestamp 1649977179
transform 1 0 25576 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0638_
timestamp 1649977179
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0639_
timestamp 1649977179
transform 1 0 25300 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0640_
timestamp 1649977179
transform -1 0 22816 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0641_
timestamp 1649977179
transform -1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0642_
timestamp 1649977179
transform 1 0 24748 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0643_
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _0644_
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0645_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21436 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0646_
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0647_
timestamp 1649977179
transform -1 0 12880 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1649977179
transform -1 0 29072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1649977179
transform 1 0 7544 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1649977179
transform -1 0 4692 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1649977179
transform -1 0 9292 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1649977179
transform -1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1649977179
transform -1 0 7544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1649977179
transform -1 0 6716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1649977179
transform -1 0 36800 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0658_
timestamp 1649977179
transform 1 0 37536 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1649977179
transform -1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0660_
timestamp 1649977179
transform 1 0 21896 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0661_
timestamp 1649977179
transform 1 0 29808 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0662_
timestamp 1649977179
transform -1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0663_
timestamp 1649977179
transform -1 0 40204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1649977179
transform -1 0 37904 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0665_
timestamp 1649977179
transform -1 0 31188 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0666_
timestamp 1649977179
transform 1 0 38732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0667_
timestamp 1649977179
transform -1 0 33120 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0668_
timestamp 1649977179
transform -1 0 32936 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0669_
timestamp 1649977179
transform -1 0 30084 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1649977179
transform -1 0 31280 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0671_
timestamp 1649977179
transform -1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0672_
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1649977179
transform 1 0 36248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1649977179
transform -1 0 34224 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0675_
timestamp 1649977179
transform -1 0 37628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1649977179
transform -1 0 34224 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0677_
timestamp 1649977179
transform -1 0 42780 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 1649977179
transform -1 0 44528 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0679_
timestamp 1649977179
transform -1 0 33488 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0680_
timestamp 1649977179
transform -1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1649977179
transform -1 0 33764 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1649977179
transform -1 0 31648 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0683_
timestamp 1649977179
transform -1 0 40572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0684_
timestamp 1649977179
transform -1 0 41768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1649977179
transform -1 0 39376 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0686_
timestamp 1649977179
transform -1 0 39284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0687_
timestamp 1649977179
transform -1 0 35052 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1649977179
transform 1 0 36432 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0690_
timestamp 1649977179
transform -1 0 30084 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1649977179
transform -1 0 26496 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0692_
timestamp 1649977179
transform -1 0 27508 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1649977179
transform -1 0 38548 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0695_
timestamp 1649977179
transform -1 0 40112 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0696_
timestamp 1649977179
transform -1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0697_
timestamp 1649977179
transform -1 0 39376 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0698_
timestamp 1649977179
transform 1 0 39652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0699_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28428 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0700_
timestamp 1649977179
transform 1 0 35788 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0701_
timestamp 1649977179
transform -1 0 30176 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0702_
timestamp 1649977179
transform -1 0 31556 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  _0703_
timestamp 1649977179
transform -1 0 28612 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0704_
timestamp 1649977179
transform 1 0 28980 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0705_
timestamp 1649977179
transform -1 0 30268 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1649977179
transform 1 0 39008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0707_
timestamp 1649977179
transform 1 0 3680 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1649977179
transform -1 0 4048 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0709_
timestamp 1649977179
transform -1 0 17020 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0710_
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _0711_
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1649977179
transform -1 0 27600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1649977179
transform -1 0 17756 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0714_
timestamp 1649977179
transform 1 0 19320 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1649977179
transform -1 0 5336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1649977179
transform -1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1649977179
transform -1 0 8464 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1649977179
transform -1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1649977179
transform -1 0 4692 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1649977179
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1649977179
transform -1 0 11040 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1649977179
transform -1 0 9568 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1649977179
transform -1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1649977179
transform -1 0 10396 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1649977179
transform -1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1649977179
transform -1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 1649977179
transform -1 0 10396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1649977179
transform -1 0 9752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1649977179
transform -1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1649977179
transform -1 0 17480 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1649977179
transform -1 0 21252 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1649977179
transform 1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1649977179
transform -1 0 19780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1649977179
transform -1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1649977179
transform -1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0741_
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1649977179
transform -1 0 20516 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1649977179
transform 1 0 23368 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1649977179
transform -1 0 22080 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1649977179
transform 1 0 22724 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1649977179
transform -1 0 18768 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1649977179
transform -1 0 19964 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1649977179
transform -1 0 20424 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1649977179
transform 1 0 22632 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1649977179
transform 1 0 27968 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1649977179
transform -1 0 27600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0753_
timestamp 1649977179
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1649977179
transform 1 0 28152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0755_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0756_
timestamp 1649977179
transform 1 0 7268 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0757_
timestamp 1649977179
transform 1 0 6440 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0758_
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0759_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 52256 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0760_
timestamp 1649977179
transform -1 0 53268 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0761_
timestamp 1649977179
transform -1 0 48576 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0762_
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 1649977179
transform 1 0 48852 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0764_
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0765_
timestamp 1649977179
transform 1 0 51428 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0766_
timestamp 1649977179
transform -1 0 53360 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0767_
timestamp 1649977179
transform -1 0 53268 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0768_
timestamp 1649977179
transform -1 0 51152 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0769_
timestamp 1649977179
transform 1 0 44804 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0770_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 48944 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0772_
timestamp 1649977179
transform 1 0 44436 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0773_
timestamp 1649977179
transform 1 0 47380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0774_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 48576 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0775_
timestamp 1649977179
transform 1 0 48116 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0776_
timestamp 1649977179
transform 1 0 44712 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0777_
timestamp 1649977179
transform -1 0 46828 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0778_
timestamp 1649977179
transform -1 0 43516 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0779_
timestamp 1649977179
transform 1 0 45908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0780_
timestamp 1649977179
transform 1 0 43884 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1649977179
transform 1 0 48944 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0782_
timestamp 1649977179
transform -1 0 48484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0783_
timestamp 1649977179
transform 1 0 48116 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0784_
timestamp 1649977179
transform -1 0 44528 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0785_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0786_
timestamp 1649977179
transform 1 0 45816 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0787_
timestamp 1649977179
transform 1 0 46644 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0788_
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0789_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 45080 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1649977179
transform -1 0 44988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0791_
timestamp 1649977179
transform -1 0 45632 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0792_
timestamp 1649977179
transform -1 0 50416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0793_
timestamp 1649977179
transform 1 0 47012 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0794_
timestamp 1649977179
transform 1 0 43884 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0795_
timestamp 1649977179
transform -1 0 50784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0796_
timestamp 1649977179
transform 1 0 48760 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0797_
timestamp 1649977179
transform -1 0 49496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0798_
timestamp 1649977179
transform 1 0 48116 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0799_
timestamp 1649977179
transform 1 0 43976 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0800_
timestamp 1649977179
transform 1 0 50784 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0801_
timestamp 1649977179
transform 1 0 51152 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0803_
timestamp 1649977179
transform -1 0 52348 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0804_
timestamp 1649977179
transform -1 0 54096 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0805_
timestamp 1649977179
transform 1 0 51704 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0806_
timestamp 1649977179
transform 1 0 51520 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0807_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 53268 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0808_
timestamp 1649977179
transform 1 0 54004 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0809_
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1649977179
transform -1 0 51060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1649977179
transform 1 0 51428 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0812_
timestamp 1649977179
transform -1 0 51336 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0813_
timestamp 1649977179
transform -1 0 57408 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0814_
timestamp 1649977179
transform 1 0 50416 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0815_
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0816_
timestamp 1649977179
transform 1 0 54096 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0817_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 54280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0818_
timestamp 1649977179
transform 1 0 53636 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0819_
timestamp 1649977179
transform 1 0 55568 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0820_
timestamp 1649977179
transform -1 0 55200 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0821_
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0823_
timestamp 1649977179
transform 1 0 47932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0824_
timestamp 1649977179
transform -1 0 55568 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0825_
timestamp 1649977179
transform 1 0 56120 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0826_
timestamp 1649977179
transform 1 0 47288 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0827_
timestamp 1649977179
transform -1 0 43332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0828_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0829_
timestamp 1649977179
transform -1 0 44712 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0830_
timestamp 1649977179
transform -1 0 50784 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0831_
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0832_
timestamp 1649977179
transform 1 0 25300 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0833_
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0834_
timestamp 1649977179
transform 1 0 40756 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0835_
timestamp 1649977179
transform 1 0 37168 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0836_
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0837_
timestamp 1649977179
transform 1 0 31188 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0838_
timestamp 1649977179
transform 1 0 26220 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0839_
timestamp 1649977179
transform 1 0 35144 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0840_
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_1  _0841_
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0842_
timestamp 1649977179
transform 1 0 53912 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0843_
timestamp 1649977179
transform -1 0 54464 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0844_
timestamp 1649977179
transform -1 0 50692 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0845_
timestamp 1649977179
transform -1 0 49680 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0846_
timestamp 1649977179
transform -1 0 52164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0847_
timestamp 1649977179
transform 1 0 51060 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0848_
timestamp 1649977179
transform 1 0 51428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0849_
timestamp 1649977179
transform -1 0 53544 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0850_
timestamp 1649977179
transform -1 0 53544 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0851_
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0852_
timestamp 1649977179
transform -1 0 48024 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0853_
timestamp 1649977179
transform 1 0 48208 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0854_
timestamp 1649977179
transform 1 0 44252 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0855_
timestamp 1649977179
transform -1 0 49588 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0856_
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0857_
timestamp 1649977179
transform -1 0 48944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0858_
timestamp 1649977179
transform 1 0 48024 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0859_
timestamp 1649977179
transform 1 0 51060 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0860_
timestamp 1649977179
transform -1 0 50692 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0861_
timestamp 1649977179
transform 1 0 50692 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0862_
timestamp 1649977179
transform -1 0 53912 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0863_
timestamp 1649977179
transform 1 0 53728 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0864_
timestamp 1649977179
transform 1 0 54004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0865_
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0866_
timestamp 1649977179
transform 1 0 51704 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0867_
timestamp 1649977179
transform -1 0 51888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0868_
timestamp 1649977179
transform 1 0 51244 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0869_
timestamp 1649977179
transform 1 0 52072 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0870_
timestamp 1649977179
transform -1 0 53268 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0871_
timestamp 1649977179
transform 1 0 52716 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0872_
timestamp 1649977179
transform -1 0 52532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0873_
timestamp 1649977179
transform 1 0 52716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0874_
timestamp 1649977179
transform 1 0 53728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0875_
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0876_
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0877_
timestamp 1649977179
transform -1 0 51520 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0878_
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0879_
timestamp 1649977179
transform 1 0 51612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0880_
timestamp 1649977179
transform -1 0 54372 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0881_
timestamp 1649977179
transform 1 0 55384 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0882_
timestamp 1649977179
transform 1 0 53912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0883_
timestamp 1649977179
transform 1 0 53084 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0884_
timestamp 1649977179
transform 1 0 54096 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1649977179
transform -1 0 54004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1649977179
transform -1 0 53544 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0887_
timestamp 1649977179
transform 1 0 53084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0888_
timestamp 1649977179
transform 1 0 54740 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0889_
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0890_
timestamp 1649977179
transform -1 0 52716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0891_
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0892_
timestamp 1649977179
transform -1 0 49772 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0893_
timestamp 1649977179
transform 1 0 47932 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0894_
timestamp 1649977179
transform 1 0 48760 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0895_
timestamp 1649977179
transform 1 0 45356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0896_
timestamp 1649977179
transform 1 0 48484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0897_
timestamp 1649977179
transform 1 0 52808 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0898_
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0899_
timestamp 1649977179
transform -1 0 48392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0900_
timestamp 1649977179
transform 1 0 48852 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0901_
timestamp 1649977179
transform -1 0 48208 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0902_
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0903_
timestamp 1649977179
transform -1 0 45632 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0904_
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0905_
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0906_
timestamp 1649977179
transform 1 0 34408 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0907_
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0908_
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0909_
timestamp 1649977179
transform 1 0 40848 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0910_
timestamp 1649977179
transform 1 0 34868 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0911_
timestamp 1649977179
transform 1 0 30452 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0912_
timestamp 1649977179
transform 1 0 27692 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0913_
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0914_
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0915_
timestamp 1649977179
transform 1 0 5060 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0916_
timestamp 1649977179
transform -1 0 6256 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0917_
timestamp 1649977179
transform 1 0 4968 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0918_
timestamp 1649977179
transform 1 0 6164 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0919_
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0920_
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0922_
timestamp 1649977179
transform 1 0 19964 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0923_
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0924_
timestamp 1649977179
transform -1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1649977179
transform -1 0 38640 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0926_
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0927_
timestamp 1649977179
transform 1 0 22172 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0928_
timestamp 1649977179
transform -1 0 27140 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0929_
timestamp 1649977179
transform 1 0 27232 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0930_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0931_
timestamp 1649977179
transform 1 0 24564 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1649977179
transform 1 0 21620 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0933_
timestamp 1649977179
transform 1 0 23276 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0934_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0935_
timestamp 1649977179
transform 1 0 24472 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0936_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25668 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _0937_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0938_
timestamp 1649977179
transform 1 0 27968 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0939_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27692 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0940_
timestamp 1649977179
transform -1 0 29072 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0941_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27968 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0942_
timestamp 1649977179
transform 1 0 29256 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0943_
timestamp 1649977179
transform 1 0 28152 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _0944_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0945_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 26404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0946_
timestamp 1649977179
transform 1 0 25668 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0947_
timestamp 1649977179
transform 1 0 4876 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0948_
timestamp 1649977179
transform 1 0 17664 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0949_
timestamp 1649977179
transform 1 0 27048 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0950_
timestamp 1649977179
transform 1 0 19688 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_1  _0951_
timestamp 1649977179
transform -1 0 42964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0952_
timestamp 1649977179
transform 1 0 38732 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0953_
timestamp 1649977179
transform -1 0 31740 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0954_
timestamp 1649977179
transform 1 0 31004 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0955_
timestamp 1649977179
transform 1 0 35972 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0956_
timestamp 1649977179
transform -1 0 41860 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0957_
timestamp 1649977179
transform -1 0 37812 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0958_
timestamp 1649977179
transform -1 0 31648 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0959_
timestamp 1649977179
transform -1 0 31004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0960_
timestamp 1649977179
transform 1 0 35328 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0961_
timestamp 1649977179
transform -1 0 40388 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0962_
timestamp 1649977179
transform -1 0 39192 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0963_
timestamp 1649977179
transform -1 0 31280 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0964_
timestamp 1649977179
transform -1 0 31648 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0965_
timestamp 1649977179
transform 1 0 30268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0966_
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0967_
timestamp 1649977179
transform -1 0 34960 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0968_
timestamp 1649977179
transform 1 0 33396 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0969_
timestamp 1649977179
transform 1 0 33488 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1649977179
transform -1 0 31004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0971_
timestamp 1649977179
transform 1 0 29992 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0972_
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0973_
timestamp 1649977179
transform 1 0 31004 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0974_
timestamp 1649977179
transform -1 0 41584 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0975_
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0976_
timestamp 1649977179
transform -1 0 28796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0977_
timestamp 1649977179
transform 1 0 28152 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0978_
timestamp 1649977179
transform 1 0 32384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0979_
timestamp 1649977179
transform -1 0 33028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0980_
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0981_
timestamp 1649977179
transform -1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0982_
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0983_
timestamp 1649977179
transform 1 0 30452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0984_
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0985_
timestamp 1649977179
transform 1 0 27876 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0986_
timestamp 1649977179
transform -1 0 27508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0987_
timestamp 1649977179
transform 1 0 26220 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1649977179
transform 1 0 31832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0989_
timestamp 1649977179
transform -1 0 43976 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0990_
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0991_
timestamp 1649977179
transform 1 0 30820 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0992_
timestamp 1649977179
transform -1 0 38548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0993_
timestamp 1649977179
transform -1 0 33580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0994_
timestamp 1649977179
transform 1 0 30544 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1649977179
transform -1 0 40112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0997_
timestamp 1649977179
transform -1 0 37996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0998_
timestamp 1649977179
transform -1 0 37904 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0999_
timestamp 1649977179
transform -1 0 41768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1000_
timestamp 1649977179
transform -1 0 38640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1001_
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1002_
timestamp 1649977179
transform -1 0 41308 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1003_
timestamp 1649977179
transform -1 0 44436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1649977179
transform 1 0 42412 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1649977179
transform 1 0 43240 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1006_
timestamp 1649977179
transform 1 0 42320 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1007_
timestamp 1649977179
transform 1 0 41032 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1008_
timestamp 1649977179
transform -1 0 42044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1009_
timestamp 1649977179
transform -1 0 43240 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1010_
timestamp 1649977179
transform -1 0 44252 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1011_
timestamp 1649977179
transform -1 0 40204 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1012_
timestamp 1649977179
transform 1 0 38180 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1013_
timestamp 1649977179
transform -1 0 37812 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1014_
timestamp 1649977179
transform -1 0 40480 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1015_
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1016_
timestamp 1649977179
transform 1 0 5704 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1017_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1018_
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _1019_
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1020_
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1021_
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1022_
timestamp 1649977179
transform 1 0 12144 0 -1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _1023_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1024_
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_2  _1025_
timestamp 1649977179
transform -1 0 44712 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1026_
timestamp 1649977179
transform -1 0 40388 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1027_
timestamp 1649977179
transform -1 0 35512 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1028_
timestamp 1649977179
transform 1 0 27784 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1029_
timestamp 1649977179
transform 1 0 28428 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1030_
timestamp 1649977179
transform -1 0 45724 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1031_
timestamp 1649977179
transform -1 0 41032 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1032_
timestamp 1649977179
transform -1 0 36892 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1033_
timestamp 1649977179
transform 1 0 27968 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1034_
timestamp 1649977179
transform 1 0 30452 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1035_
timestamp 1649977179
transform -1 0 32844 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1036_
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1037_
timestamp 1649977179
transform -1 0 29440 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1038_
timestamp 1649977179
transform -1 0 30084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1039_
timestamp 1649977179
transform 1 0 28704 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1040_
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 1649977179
transform 1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1042_
timestamp 1649977179
transform 1 0 30268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1043_
timestamp 1649977179
transform 1 0 28520 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1044_
timestamp 1649977179
transform -1 0 27600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1045_
timestamp 1649977179
transform 1 0 28152 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1046_
timestamp 1649977179
transform -1 0 29440 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1047_
timestamp 1649977179
transform 1 0 28428 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1048_
timestamp 1649977179
transform -1 0 28612 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1049_
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1050_
timestamp 1649977179
transform 1 0 30820 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1649977179
transform 1 0 33396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1052_
timestamp 1649977179
transform -1 0 34224 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1053_
timestamp 1649977179
transform 1 0 34224 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1054_
timestamp 1649977179
transform -1 0 39192 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1055_
timestamp 1649977179
transform 1 0 31372 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1056_
timestamp 1649977179
transform -1 0 31832 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1057_
timestamp 1649977179
transform 1 0 30912 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1058_
timestamp 1649977179
transform 1 0 38548 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1059_
timestamp 1649977179
transform -1 0 37812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1060_
timestamp 1649977179
transform 1 0 38272 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1061_
timestamp 1649977179
transform -1 0 39376 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1062_
timestamp 1649977179
transform -1 0 36800 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1063_
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1064_
timestamp 1649977179
transform -1 0 37904 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1065_
timestamp 1649977179
transform 1 0 40664 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1066_
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1649977179
transform -1 0 41492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1068_
timestamp 1649977179
transform -1 0 40664 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1070_
timestamp 1649977179
transform 1 0 41216 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1071_
timestamp 1649977179
transform -1 0 42780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1072_
timestamp 1649977179
transform 1 0 39928 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1073_
timestamp 1649977179
transform -1 0 44528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1074_
timestamp 1649977179
transform -1 0 46920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1075_
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1076_
timestamp 1649977179
transform 1 0 46920 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1077_
timestamp 1649977179
transform 1 0 46184 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1078_
timestamp 1649977179
transform -1 0 45816 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1079_
timestamp 1649977179
transform 1 0 45816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1080_
timestamp 1649977179
transform 1 0 46000 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1081_
timestamp 1649977179
transform -1 0 45632 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1082_
timestamp 1649977179
transform 1 0 30268 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1083_
timestamp 1649977179
transform 1 0 30360 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1084_
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1085_
timestamp 1649977179
transform 1 0 39652 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1086_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1087_
timestamp 1649977179
transform 1 0 21896 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1088_
timestamp 1649977179
transform 1 0 20148 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1089_
timestamp 1649977179
transform 1 0 27324 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1090_
timestamp 1649977179
transform 1 0 27876 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1091_
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1092_
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1093_
timestamp 1649977179
transform 1 0 25300 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1094_
timestamp 1649977179
transform 1 0 27324 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1095_
timestamp 1649977179
transform 1 0 28888 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1096_
timestamp 1649977179
transform 1 0 17388 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1097_
timestamp 1649977179
transform -1 0 18124 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1098_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1099_
timestamp 1649977179
transform 1 0 17940 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1100_
timestamp 1649977179
transform -1 0 5428 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1101_
timestamp 1649977179
transform 1 0 26312 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1103_
timestamp 1649977179
transform 1 0 25392 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1104_
timestamp 1649977179
transform 1 0 25852 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1105_
timestamp 1649977179
transform -1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1106_
timestamp 1649977179
transform -1 0 33396 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1107_
timestamp 1649977179
transform 1 0 23828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1108_
timestamp 1649977179
transform -1 0 23000 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1109_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1110_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27048 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1111_
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1112_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23920 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1113_
timestamp 1649977179
transform -1 0 19964 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__or3_1  _1114_
timestamp 1649977179
transform 1 0 25668 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1115_
timestamp 1649977179
transform 1 0 25760 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1116_
timestamp 1649977179
transform -1 0 25392 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1117_
timestamp 1649977179
transform -1 0 25668 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1118__29
timestamp 1649977179
transform -1 0 5888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119__30
timestamp 1649977179
transform 1 0 7176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1120_
timestamp 1649977179
transform 1 0 4324 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121__31
timestamp 1649977179
transform 1 0 4784 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122__32
timestamp 1649977179
transform -1 0 4876 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1123__33
timestamp 1649977179
transform -1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1124__34
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125__35
timestamp 1649977179
transform 1 0 7912 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1126_
timestamp 1649977179
transform 1 0 10580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127__36
timestamp 1649977179
transform 1 0 11684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128__37
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129__38
timestamp 1649977179
transform -1 0 16100 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1130__39
timestamp 1649977179
transform -1 0 14260 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131__40
timestamp 1649977179
transform -1 0 16192 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1132_
timestamp 1649977179
transform 1 0 12696 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1133_
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1134__41
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1135__42
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1136__43
timestamp 1649977179
transform 1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1137_
timestamp 1649977179
transform 1 0 2944 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1138_
timestamp 1649977179
transform 1 0 1932 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1139__44
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1140_
timestamp 1649977179
transform 1 0 1932 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1141__45
timestamp 1649977179
transform -1 0 9384 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1142_
timestamp 1649977179
transform 1 0 1932 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1143_
timestamp 1649977179
transform -1 0 35788 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1649977179
transform -1 0 39744 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1649977179
transform -1 0 24656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1649977179
transform -1 0 32384 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1649977179
transform -1 0 40848 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1649977179
transform -1 0 42688 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1149_
timestamp 1649977179
transform -1 0 34500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1150_
timestamp 1649977179
transform -1 0 33580 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1649977179
transform 1 0 30452 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1649977179
transform -1 0 29808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1153_
timestamp 1649977179
transform -1 0 35512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1155_
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1156_
timestamp 1649977179
transform 1 0 36984 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1649977179
transform 1 0 40296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1158_
timestamp 1649977179
transform -1 0 34960 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1159_
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1649977179
transform -1 0 35604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1161_
timestamp 1649977179
transform 1 0 22264 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1649977179
transform 1 0 41124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1163_
timestamp 1649977179
transform 1 0 19320 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1164_
timestamp 1649977179
transform 1 0 20976 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1649977179
transform -1 0 40480 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1166_
timestamp 1649977179
transform 1 0 19320 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1167_
timestamp 1649977179
transform -1 0 36524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1649977179
transform -1 0 34132 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1169_
timestamp 1649977179
transform 1 0 16928 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1649977179
transform -1 0 31280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1171_
timestamp 1649977179
transform 1 0 12052 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1649977179
transform -1 0 28520 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1649977179
transform 1 0 38088 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1174_
timestamp 1649977179
transform 1 0 20240 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1176_
timestamp 1649977179
transform 1 0 17848 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1177_
timestamp 1649977179
transform -1 0 36156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1178_
timestamp 1649977179
transform 1 0 15272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1179__46
timestamp 1649977179
transform -1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1180__47
timestamp 1649977179
transform 1 0 19504 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1181_
timestamp 1649977179
transform 1 0 14168 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1182_
timestamp 1649977179
transform 1 0 14720 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1183_
timestamp 1649977179
transform 1 0 14444 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1184__48
timestamp 1649977179
transform 1 0 16744 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1185_
timestamp 1649977179
transform -1 0 7820 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1186__49
timestamp 1649977179
transform 1 0 15364 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1187_
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1188__50
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1189_
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1190_
timestamp 1649977179
transform -1 0 16192 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1191_
timestamp 1649977179
transform -1 0 12512 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1192__51
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1193_
timestamp 1649977179
transform -1 0 14904 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1194__52
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1195_
timestamp 1649977179
transform -1 0 15272 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1196__53
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1197_
timestamp 1649977179
transform 1 0 9752 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1198__54
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1199__55
timestamp 1649977179
transform -1 0 10948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1200_
timestamp 1649977179
transform 1 0 7636 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1201_
timestamp 1649977179
transform 1 0 14444 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1202__56
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1203_
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1204__57
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1205_
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1206__58
timestamp 1649977179
transform -1 0 11868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1207_
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1208__59
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1209_
timestamp 1649977179
transform 1 0 20884 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1210__60
timestamp 1649977179
transform -1 0 18584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1211_
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1212_
timestamp 1649977179
transform 1 0 21988 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _1213_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1214__61
timestamp 1649977179
transform -1 0 14996 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1215_
timestamp 1649977179
transform 1 0 18124 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1216__62
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1217_
timestamp 1649977179
transform 1 0 14536 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1218__63
timestamp 1649977179
transform -1 0 17480 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1219_
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1220__64
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1221__65
timestamp 1649977179
transform 1 0 17848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1222_
timestamp 1649977179
transform 1 0 19412 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1223__3
timestamp 1649977179
transform 1 0 25392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1224_
timestamp 1649977179
transform 1 0 17296 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1225__4
timestamp 1649977179
transform -1 0 26864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1226_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1227__5
timestamp 1649977179
transform -1 0 25576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1228_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 1649977179
transform -1 0 5888 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1230_
timestamp 1649977179
transform -1 0 8464 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1231_
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1232_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1233_
timestamp 1649977179
transform 1 0 6716 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1234_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1235_
timestamp 1649977179
transform 1 0 6532 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1236_
timestamp 1649977179
transform -1 0 3220 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1237_
timestamp 1649977179
transform 1 0 9200 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1238_
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 1649977179
transform 1 0 8924 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1240_
timestamp 1649977179
transform 1 0 9200 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1241_
timestamp 1649977179
transform 1 0 6716 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1242_
timestamp 1649977179
transform 1 0 13800 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1243_
timestamp 1649977179
transform 1 0 11776 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 1649977179
transform 1 0 18032 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1245_
timestamp 1649977179
transform -1 0 13524 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1246_
timestamp 1649977179
transform 1 0 22080 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1247_
timestamp 1649977179
transform -1 0 15916 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1248_
timestamp 1649977179
transform 1 0 19320 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1249_
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1250_
timestamp 1649977179
transform 1 0 27232 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1251_
timestamp 1649977179
transform -1 0 15916 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1252_
timestamp 1649977179
transform 1 0 22448 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1253_
timestamp 1649977179
transform 1 0 12144 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1254_
timestamp 1649977179
transform -1 0 11040 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1255_
timestamp 1649977179
transform -1 0 3680 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1256_
timestamp 1649977179
transform -1 0 11040 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1257_
timestamp 1649977179
transform 1 0 3864 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1258_
timestamp 1649977179
transform -1 0 11040 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1259_
timestamp 1649977179
transform 1 0 3496 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1260_
timestamp 1649977179
transform -1 0 12236 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1261_
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1262_
timestamp 1649977179
transform -1 0 50508 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1263_
timestamp 1649977179
transform 1 0 45356 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1264_
timestamp 1649977179
transform 1 0 48944 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1265_
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1266_
timestamp 1649977179
transform 1 0 44436 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1267_
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1268_
timestamp 1649977179
transform -1 0 49036 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1269_
timestamp 1649977179
transform -1 0 52164 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1270_
timestamp 1649977179
transform 1 0 51612 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1271_
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1272_
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1273_
timestamp 1649977179
transform -1 0 56948 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1274_
timestamp 1649977179
transform 1 0 56304 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1275_
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1276_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 44252 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1277_
timestamp 1649977179
transform 1 0 49404 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1278_
timestamp 1649977179
transform -1 0 36984 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1279_
timestamp 1649977179
transform -1 0 39100 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1280_
timestamp 1649977179
transform 1 0 19872 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1281_
timestamp 1649977179
transform 1 0 22080 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1282_
timestamp 1649977179
transform 1 0 30544 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1283_
timestamp 1649977179
transform 1 0 27784 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1284_
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 1649977179
transform 1 0 36340 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 1649977179
transform 1 0 29348 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 1649977179
transform -1 0 38088 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1288_
timestamp 1649977179
transform 1 0 31096 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1289_
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1290_
timestamp 1649977179
transform 1 0 29808 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1291_
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1292_
timestamp 1649977179
transform 1 0 23276 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1293_
timestamp 1649977179
transform -1 0 26036 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1294_
timestamp 1649977179
transform -1 0 35880 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1295_
timestamp 1649977179
transform 1 0 33672 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1296_
timestamp 1649977179
transform -1 0 36800 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1297_
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1298_
timestamp 1649977179
transform 1 0 45264 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1299_
timestamp 1649977179
transform 1 0 48392 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1300_
timestamp 1649977179
transform 1 0 51704 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1301_
timestamp 1649977179
transform 1 0 55384 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1302_
timestamp 1649977179
transform 1 0 51704 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1303_
timestamp 1649977179
transform 1 0 54280 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1304_
timestamp 1649977179
transform 1 0 56304 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1305_
timestamp 1649977179
transform -1 0 50876 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1306_
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1307_
timestamp 1649977179
transform -1 0 55660 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1308_
timestamp 1649977179
transform -1 0 58236 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1309_
timestamp 1649977179
transform -1 0 57132 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1310_
timestamp 1649977179
transform 1 0 54280 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1311_
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1312_
timestamp 1649977179
transform 1 0 44712 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 1649977179
transform 1 0 48852 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 1649977179
transform 1 0 41584 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1315_
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1316_
timestamp 1649977179
transform 1 0 32200 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1317_
timestamp 1649977179
transform 1 0 31004 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1318_
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1319_
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1320_
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1321_
timestamp 1649977179
transform 1 0 39192 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1322_
timestamp 1649977179
transform 1 0 36708 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1323_
timestamp 1649977179
transform 1 0 37996 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1324_
timestamp 1649977179
transform 1 0 33580 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1325_
timestamp 1649977179
transform 1 0 32384 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1326_
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1327_
timestamp 1649977179
transform 1 0 29900 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1328_
timestamp 1649977179
transform 1 0 26312 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1329_
timestamp 1649977179
transform 1 0 26496 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1330_
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1331_
timestamp 1649977179
transform 1 0 37352 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1332_
timestamp 1649977179
transform 1 0 37996 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1333_
timestamp 1649977179
transform -1 0 41676 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1334_
timestamp 1649977179
transform 1 0 6992 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1335_
timestamp 1649977179
transform -1 0 4140 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1336_
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1338_
timestamp 1649977179
transform -1 0 58144 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1339_
timestamp 1649977179
transform -1 0 57408 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1340_
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1341_
timestamp 1649977179
transform 1 0 18400 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1342_
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1343_
timestamp 1649977179
transform 1 0 35880 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1344_
timestamp 1649977179
transform 1 0 19412 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1345_
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1346_
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1347_
timestamp 1649977179
transform -1 0 5612 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1348_
timestamp 1649977179
transform -1 0 3312 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1349_
timestamp 1649977179
transform 1 0 15732 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1350_
timestamp 1649977179
transform -1 0 20700 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1351_
timestamp 1649977179
transform 1 0 26864 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1352_
timestamp 1649977179
transform 1 0 24656 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1353_
timestamp 1649977179
transform 1 0 16192 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1354_
timestamp 1649977179
transform -1 0 21068 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1355_
timestamp 1649977179
transform -1 0 39192 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1356_
timestamp 1649977179
transform 1 0 33580 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1357_
timestamp 1649977179
transform 1 0 33764 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1358_
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1359_
timestamp 1649977179
transform 1 0 33856 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1360_
timestamp 1649977179
transform 1 0 35052 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1361_
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1362_
timestamp 1649977179
transform 1 0 33672 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1363_
timestamp 1649977179
transform 1 0 32660 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1364_
timestamp 1649977179
transform 1 0 34868 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1365_
timestamp 1649977179
transform 1 0 37260 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1366_
timestamp 1649977179
transform 1 0 38824 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1367_
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1368_
timestamp 1649977179
transform -1 0 43516 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1369_
timestamp 1649977179
transform -1 0 37536 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1370_
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1371_
timestamp 1649977179
transform -1 0 19320 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1372_
timestamp 1649977179
transform 1 0 6532 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1373_
timestamp 1649977179
transform -1 0 19044 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1374_
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1375_
timestamp 1649977179
transform -1 0 21160 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1376_
timestamp 1649977179
transform 1 0 6992 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1377_
timestamp 1649977179
transform -1 0 8280 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1378_
timestamp 1649977179
transform -1 0 13616 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1379_
timestamp 1649977179
transform -1 0 13432 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1380_
timestamp 1649977179
transform 1 0 9568 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1381_
timestamp 1649977179
transform -1 0 13432 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1382_
timestamp 1649977179
transform 1 0 11960 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1383_
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1384_
timestamp 1649977179
transform -1 0 13340 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1385_
timestamp 1649977179
transform -1 0 13248 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1386_
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1387_
timestamp 1649977179
transform -1 0 17020 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1388_
timestamp 1649977179
transform 1 0 9384 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1389_
timestamp 1649977179
transform -1 0 16100 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1390_
timestamp 1649977179
transform 1 0 22080 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1391_
timestamp 1649977179
transform 1 0 32384 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1392_
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1393_
timestamp 1649977179
transform -1 0 36524 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1394_
timestamp 1649977179
transform 1 0 32384 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1395_
timestamp 1649977179
transform -1 0 35144 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1396_
timestamp 1649977179
transform 1 0 35328 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1397_
timestamp 1649977179
transform 1 0 33304 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1398_
timestamp 1649977179
transform -1 0 40112 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1399_
timestamp 1649977179
transform -1 0 38824 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1400_
timestamp 1649977179
transform -1 0 43056 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1401_
timestamp 1649977179
transform -1 0 42780 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1402_
timestamp 1649977179
transform -1 0 43332 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1403_
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1404_
timestamp 1649977179
transform 1 0 42320 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1405_
timestamp 1649977179
transform -1 0 35328 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1406_
timestamp 1649977179
transform 1 0 40112 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1407_
timestamp 1649977179
transform -1 0 16100 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1408_
timestamp 1649977179
transform 1 0 23460 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1409_
timestamp 1649977179
transform -1 0 20332 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1410_
timestamp 1649977179
transform 1 0 22080 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1411_
timestamp 1649977179
transform 1 0 14352 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1412_
timestamp 1649977179
transform -1 0 26220 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1413_
timestamp 1649977179
transform 1 0 22172 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1414_
timestamp 1649977179
transform -1 0 17940 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1415_
timestamp 1649977179
transform 1 0 24380 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1416_
timestamp 1649977179
transform 1 0 15916 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1417_
timestamp 1649977179
transform 1 0 23276 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1418_
timestamp 1649977179
transform 1 0 16008 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1419_
timestamp 1649977179
transform 1 0 22080 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1420_
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1421_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1422_
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1423_
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1424_
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1425_
timestamp 1649977179
transform 1 0 24380 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1426_
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1427_
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1428_
timestamp 1649977179
transform -1 0 20792 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1429_
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1430_
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1431_
timestamp 1649977179
transform -1 0 39100 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1432_
timestamp 1649977179
transform -1 0 29072 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1433_
timestamp 1649977179
transform -1 0 24932 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1434_
timestamp 1649977179
transform 1 0 25392 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1435_
timestamp 1649977179
transform 1 0 25944 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  _1436_
timestamp 1649977179
transform 1 0 33304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1437_
timestamp 1649977179
transform 1 0 41400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1438_
timestamp 1649977179
transform 1 0 43700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1439_
timestamp 1649977179
transform -1 0 57408 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1440_
timestamp 1649977179
transform 1 0 37720 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1649977179
transform -1 0 47104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1442_
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1649977179
transform -1 0 47656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1444_
timestamp 1649977179
transform -1 0 4600 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1649977179
transform 1 0 2208 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1447_
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1448_
timestamp 1649977179
transform 1 0 2852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1649977179
transform -1 0 40112 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1451_
timestamp 1649977179
transform -1 0 25024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1452_
timestamp 1649977179
transform 1 0 13064 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1649977179
transform 1 0 17480 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1454_
timestamp 1649977179
transform 1 0 38088 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1455_
timestamp 1649977179
transform -1 0 49588 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1649977179
transform -1 0 48944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1649977179
transform 1 0 19596 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1458_
timestamp 1649977179
transform 1 0 2208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1459_
timestamp 1649977179
transform -1 0 46092 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1460_
timestamp 1649977179
transform -1 0 32568 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1649977179
transform -1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1462_
timestamp 1649977179
transform -1 0 2300 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1649977179
transform 1 0 22724 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0323_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6992 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0324_
timestamp 1649977179
transform 1 0 13892 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0325_
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0326_
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0332_
timestamp 1649977179
transform 1 0 18952 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0333_
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0334_
timestamp 1649977179
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0335_
timestamp 1649977179
transform 1 0 18952 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0336_
timestamp 1649977179
transform 1 0 24656 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0337_
timestamp 1649977179
transform 1 0 24932 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0338_
timestamp 1649977179
transform 1 0 24472 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0339_
timestamp 1649977179
transform -1 0 10488 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0340_
timestamp 1649977179
transform 1 0 12328 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0341_
timestamp 1649977179
transform 1 0 7820 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0348_
timestamp 1649977179
transform 1 0 4416 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_master
timestamp 1649977179
transform 1 0 19596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_w0.cclk_I
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0323_
timestamp 1649977179
transform -1 0 5888 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0324_
timestamp 1649977179
transform -1 0 12236 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0325_
timestamp 1649977179
transform -1 0 11408 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0326_
timestamp 1649977179
transform -1 0 8832 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0332_
timestamp 1649977179
transform -1 0 16468 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0333_
timestamp 1649977179
transform -1 0 12236 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0334_
timestamp 1649977179
transform -1 0 13616 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0335_
timestamp 1649977179
transform -1 0 16192 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0336_
timestamp 1649977179
transform -1 0 21712 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0337_
timestamp 1649977179
transform 1 0 22080 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0338_
timestamp 1649977179
transform -1 0 22632 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0339_
timestamp 1649977179
transform -1 0 6256 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0340_
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0341_
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0348_
timestamp 1649977179
transform -1 0 3312 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0323_
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0324_
timestamp 1649977179
transform 1 0 15640 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0325_
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0326_
timestamp 1649977179
transform -1 0 11040 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0332_
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0333_
timestamp 1649977179
transform -1 0 11040 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0334_
timestamp 1649977179
transform 1 0 14352 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0335_
timestamp 1649977179
transform 1 0 14352 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0336_
timestamp 1649977179
transform 1 0 26036 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0337_
timestamp 1649977179
transform 1 0 22172 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0338_
timestamp 1649977179
transform 1 0 22080 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0339_
timestamp 1649977179
transform 1 0 9384 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0340_
timestamp 1649977179
transform -1 0 11040 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0341_
timestamp 1649977179
transform -1 0 5980 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0348_
timestamp 1649977179
transform 1 0 6624 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk_master
timestamp 1649977179
transform -1 0 11408 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_w0.cclk_I
timestamp 1649977179
transform 1 0 35052 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk_master
timestamp 1649977179
transform -1 0 12236 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_w0.cclk_I
timestamp 1649977179
transform 1 0 39008 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk_master
timestamp 1649977179
transform 1 0 28612 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_w0.cclk_I
timestamp 1649977179
transform -1 0 35604 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk_master
timestamp 1649977179
transform 1 0 28612 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_w0.cclk_I
timestamp 1649977179
transform 1 0 39008 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 43240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 57408 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform -1 0 58236 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 24380 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1649977179
transform -1 0 53452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 28428 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform -1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  net99_2
timestamp 1649977179
transform -1 0 34040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1649977179
transform 1 0 33580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1649977179
transform -1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1649977179
transform 1 0 43240 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output15
timestamp 1649977179
transform 1 0 38732 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1649977179
transform 1 0 48392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1649977179
transform 1 0 19228 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1649977179
transform 1 0 4600 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1649977179
transform 1 0 57868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1649977179
transform -1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1649977179
transform -1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1649977179
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1649977179
transform 1 0 48392 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1649977179
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1649977179
transform -1 0 14628 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1649977179
transform 1 0 38732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform 1 0 52900 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform 1 0 57868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform -1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform 1 0 33580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform 1 0 2760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform -1 0 9476 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater39
timestamp 1649977179
transform 1 0 54280 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater40
timestamp 1649977179
transform -1 0 54832 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater41
timestamp 1649977179
transform 1 0 52808 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater42
timestamp 1649977179
transform 1 0 51060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater43
timestamp 1649977179
transform 1 0 50600 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater44
timestamp 1649977179
transform -1 0 52900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater45
timestamp 1649977179
transform -1 0 48392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater46
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater47
timestamp 1649977179
transform -1 0 50140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater48
timestamp 1649977179
transform -1 0 49496 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater49
timestamp 1649977179
transform -1 0 55660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater50
timestamp 1649977179
transform -1 0 52072 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater51
timestamp 1649977179
transform -1 0 43884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater52
timestamp 1649977179
transform -1 0 54740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater53
timestamp 1649977179
transform 1 0 51336 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater54
timestamp 1649977179
transform -1 0 51060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater55
timestamp 1649977179
transform -1 0 50416 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater56
timestamp 1649977179
transform -1 0 50416 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater57
timestamp 1649977179
transform -1 0 41952 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater58
timestamp 1649977179
transform 1 0 39008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater59
timestamp 1649977179
transform -1 0 30636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater60
timestamp 1649977179
transform -1 0 29256 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater61
timestamp 1649977179
transform 1 0 26220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater62
timestamp 1649977179
transform -1 0 16652 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater63
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater64
timestamp 1649977179
transform -1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater65
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater66
timestamp 1649977179
transform 1 0 19596 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater67
timestamp 1649977179
transform -1 0 37628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater68
timestamp 1649977179
transform -1 0 33856 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater69
timestamp 1649977179
transform 1 0 27324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater70
timestamp 1649977179
transform -1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater71
timestamp 1649977179
transform 1 0 29532 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater72
timestamp 1649977179
transform -1 0 32844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater73
timestamp 1649977179
transform 1 0 31372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater74
timestamp 1649977179
transform 1 0 31924 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater75
timestamp 1649977179
transform 1 0 35420 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater76
timestamp 1649977179
transform -1 0 35236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater77
timestamp 1649977179
transform -1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater78
timestamp 1649977179
transform 1 0 25576 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater79
timestamp 1649977179
transform -1 0 19504 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater80
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater81
timestamp 1649977179
transform 1 0 13248 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater82
timestamp 1649977179
transform 1 0 4324 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater83
timestamp 1649977179
transform 1 0 12880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater84
timestamp 1649977179
transform -1 0 18124 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater85
timestamp 1649977179
transform -1 0 43332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater86
timestamp 1649977179
transform -1 0 43332 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater87
timestamp 1649977179
transform -1 0 41860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater88
timestamp 1649977179
transform -1 0 40296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater89
timestamp 1649977179
transform 1 0 40296 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater90
timestamp 1649977179
transform -1 0 41676 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater91
timestamp 1649977179
transform -1 0 42320 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater92
timestamp 1649977179
transform -1 0 38364 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater93
timestamp 1649977179
transform -1 0 43792 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater94
timestamp 1649977179
transform -1 0 41952 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater95
timestamp 1649977179
transform -1 0 6624 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater96
timestamp 1649977179
transform -1 0 6624 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater97
timestamp 1649977179
transform -1 0 7360 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater98
timestamp 1649977179
transform -1 0 8372 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater99
timestamp 1649977179
transform -1 0 8372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater100
timestamp 1649977179
transform -1 0 8464 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater101
timestamp 1649977179
transform -1 0 10396 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater102
timestamp 1649977179
transform -1 0 13340 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater103
timestamp 1649977179
transform 1 0 14720 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater104
timestamp 1649977179
transform -1 0 15916 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater105
timestamp 1649977179
transform -1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater106
timestamp 1649977179
transform -1 0 20516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater107
timestamp 1649977179
transform -1 0 22540 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater108
timestamp 1649977179
transform 1 0 24748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater109
timestamp 1649977179
transform -1 0 23736 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater110
timestamp 1649977179
transform -1 0 25116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater111
timestamp 1649977179
transform -1 0 37536 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater112
timestamp 1649977179
transform -1 0 38180 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater113
timestamp 1649977179
transform -1 0 35420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater114
timestamp 1649977179
transform -1 0 35880 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater115
timestamp 1649977179
transform -1 0 36340 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater116
timestamp 1649977179
transform -1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater117
timestamp 1649977179
transform -1 0 40572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater118
timestamp 1649977179
transform 1 0 40480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater119
timestamp 1649977179
transform -1 0 38364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater120
timestamp 1649977179
transform -1 0 38180 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater121
timestamp 1649977179
transform 1 0 36248 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater122
timestamp 1649977179
transform -1 0 42688 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater123
timestamp 1649977179
transform 1 0 44068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater124
timestamp 1649977179
transform -1 0 42688 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater125
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater126
timestamp 1649977179
transform 1 0 53084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater127
timestamp 1649977179
transform 1 0 50048 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater128
timestamp 1649977179
transform 1 0 45356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater129
timestamp 1649977179
transform 1 0 42596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater130
timestamp 1649977179
transform 1 0 38272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater131
timestamp 1649977179
transform 1 0 36340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater132
timestamp 1649977179
transform -1 0 38180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater133
timestamp 1649977179
transform 1 0 34776 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater134
timestamp 1649977179
transform 1 0 47932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater135
timestamp 1649977179
transform -1 0 44528 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater136
timestamp 1649977179
transform -1 0 44528 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater137
timestamp 1649977179
transform -1 0 57960 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater138
timestamp 1649977179
transform 1 0 56580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater139
timestamp 1649977179
transform 1 0 50416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater140
timestamp 1649977179
transform 1 0 45080 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater141
timestamp 1649977179
transform 1 0 42320 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater142
timestamp 1649977179
transform -1 0 42688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater143
timestamp 1649977179
transform 1 0 35144 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater144
timestamp 1649977179
transform 1 0 35880 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater145
timestamp 1649977179
transform -1 0 36432 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater146
timestamp 1649977179
transform 1 0 29900 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5152 0 1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 30820 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1649977179
transform 1 0 5152 0 1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1649977179
transform 1 0 29716 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1649977179
transform 1 0 4600 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1649977179
transform -1 0 26772 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1649977179
transform -1 0 7636 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1649977179
transform 1 0 29532 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1649977179
transform -1 0 8096 0 1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1649977179
transform -1 0 8096 0 1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1649977179
transform -1 0 29072 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1649977179
transform 1 0 5152 0 1 32640
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1649977179
transform -1 0 28888 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1649977179
transform 1 0 4600 0 -1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1649977179
transform -1 0 26128 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1649977179
transform 1 0 6992 0 1 28288
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1649977179
transform -1 0 24840 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1649977179
transform 1 0 1748 0 -1 32640
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1649977179
transform -1 0 28888 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn
timestamp 1649977179
transform 1 0 36064 0 1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
timestamp 1649977179
transform -1 0 32936 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1649977179
transform 1 0 36064 0 1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1649977179
transform -1 0 30084 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1649977179
transform 1 0 35512 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1649977179
transform 1 0 34408 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1649977179
transform -1 0 38548 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1649977179
transform -1 0 39008 0 1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1649977179
transform -1 0 33856 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1649977179
transform -1 0 39008 0 1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1649977179
transform 1 0 27048 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1649977179
transform 1 0 36064 0 1 29376
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1649977179
transform 1 0 36064 0 1 32640
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1649977179
transform 1 0 16836 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1649977179
transform 1 0 35052 0 1 28288
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1649977179
transform 1 0 17112 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1649977179
transform 1 0 35144 0 -1 28288
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  w0.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  w0.ro_block_I.ro_pol.tribuf.t_buf dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  w0.ro_block_I.ro_pol_eve.tribuf.t_buf dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21344 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  w0.ro_block_Q.ro_pol.tribuf.t_buf
timestamp 1649977179
transform 1 0 5796 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  w0.ro_block_Q.ro_pol_eve.tribuf.t_buf dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43240 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
timestamp 1649977179
transform -1 0 44344 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1649977179
transform 1 0 43700 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1649977179
transform -1 0 43424 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1649977179
transform 1 0 43700 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1649977179
transform 1 0 47748 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1649977179
transform 1 0 45356 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1649977179
transform 1 0 48116 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1649977179
transform 1 0 45356 0 -1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1649977179
transform -1 0 43884 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1649977179
transform 1 0 43240 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1649977179
transform 1 0 49312 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1649977179
transform -1 0 46276 0 1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1649977179
transform -1 0 49036 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1649977179
transform -1 0 46828 0 -1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1649977179
transform -1 0 44344 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_2  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1649977179
transform -1 0 41952 0 -1 22848
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_I.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].dl.dlrtn
timestamp 1649977179
transform 1 0 40664 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[0\].t_buf.t_buf
timestamp 1649977179
transform -1 0 40572 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].dl.dlrtn
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[1\].t_buf.t_buf
timestamp 1649977179
transform -1 0 47748 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].dl.dlrtn
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[2\].t_buf.t_buf
timestamp 1649977179
transform -1 0 47104 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].dl.dlrtn
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[3\].t_buf.t_buf
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].dl.dlrtn
timestamp 1649977179
transform 1 0 42596 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[4\].t_buf.t_buf
timestamp 1649977179
transform 1 0 45172 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].dl.dlrtn
timestamp 1649977179
transform 1 0 42596 0 1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[5\].t_buf.t_buf
timestamp 1649977179
transform -1 0 43332 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].dl.dlrtn
timestamp 1649977179
transform 1 0 40664 0 -1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[6\].t_buf.t_buf
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].dl.dlrtn
timestamp 1649977179
transform 1 0 40664 0 -1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[7\].t_buf.t_buf
timestamp 1649977179
transform 1 0 37536 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].dl.dlrtn
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[8\].t_buf.t_buf
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dlrtn_1  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].dl.dlrtn
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__ebufn_8  wrapper_cell_loop\[0\].w1.fb_block_Q.gs_f.fb_gray_selector_loop\[9\].t_buf.t_buf
timestamp 1649977179
transform -1 0 45356 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  wrapper_cell_loop\[0\].w1.ro_block_I.ro_pol.tribuf.t_buf
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  wrapper_cell_loop\[0\].w1.ro_block_I.ro_pol_eve.tribuf.t_buf
timestamp 1649977179
transform -1 0 20424 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  wrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol.tribuf.t_buf
timestamp 1649977179
transform -1 0 7636 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  wrapper_cell_loop\[0\].w1.ro_block_Q.ro_pol_eve.tribuf.t_buf
timestamp 1649977179
transform 1 0 8924 0 -1 28288
box -38 -48 1234 592
<< labels >>
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 cclk_I[0]
port 0 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 cclk_I[1]
port 1 nsew signal tristate
flabel metal2 s 43166 35200 43222 36000 0 FreeSans 224 90 0 0 cclk_Q[0]
port 2 nsew signal tristate
flabel metal3 s 59200 12928 60000 13048 0 FreeSans 480 0 0 0 cclk_Q[1]
port 3 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 clk_master
port 4 nsew signal input
flabel metal2 s 38658 35200 38714 36000 0 FreeSans 224 90 0 0 clkdiv2_I[0]
port 5 nsew signal tristate
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 clkdiv2_I[1]
port 6 nsew signal tristate
flabel metal2 s 18694 35200 18750 36000 0 FreeSans 224 90 0 0 clkdiv2_Q[0]
port 7 nsew signal tristate
flabel metal3 s 59200 23128 60000 23248 0 FreeSans 480 0 0 0 clkdiv2_Q[1]
port 8 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 comp_high_I[0]
port 9 nsew signal input
flabel metal2 s 57978 35200 58034 36000 0 FreeSans 224 90 0 0 comp_high_I[1]
port 10 nsew signal input
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 comp_high_Q[0]
port 11 nsew signal input
flabel metal2 s 23846 35200 23902 36000 0 FreeSans 224 90 0 0 comp_high_Q[1]
port 12 nsew signal input
flabel metal2 s 4526 35200 4582 36000 0 FreeSans 224 90 0 0 cos_out[0]
port 13 nsew signal tristate
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 cos_out[1]
port 14 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 cos_outb[0]
port 15 nsew signal tristate
flabel metal3 s 59200 17688 60000 17808 0 FreeSans 480 0 0 0 cos_outb[1]
port 16 nsew signal tristate
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 fb1_I[0]
port 17 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 fb1_I[1]
port 18 nsew signal tristate
flabel metal2 s 48318 35200 48374 36000 0 FreeSans 224 90 0 0 fb1_Q[0]
port 19 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 fb1_Q[1]
port 20 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 fb2_I[0]
port 21 nsew signal tristate
flabel metal2 s 14186 35200 14242 36000 0 FreeSans 224 90 0 0 fb2_I[1]
port 22 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 fb2_Q[0]
port 23 nsew signal tristate
flabel metal2 s 52826 35200 52882 36000 0 FreeSans 224 90 0 0 fb2_Q[1]
port 24 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 phi1b_dig_I[0]
port 25 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 phi1b_dig_I[1]
port 26 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 phi1b_dig_Q[0]
port 27 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 phi1b_dig_Q[1]
port 28 nsew signal input
flabel metal3 s 59200 2728 60000 2848 0 FreeSans 480 0 0 0 read_out_I[0]
port 29 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 read_out_I[1]
port 30 nsew signal tristate
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 read_out_Q[0]
port 31 nsew signal tristate
flabel metal3 s 59200 33328 60000 33448 0 FreeSans 480 0 0 0 read_out_Q[1]
port 32 nsew signal tristate
flabel metal2 s 28354 35200 28410 36000 0 FreeSans 224 90 0 0 rstb
port 33 nsew signal input
flabel metal2 s 33506 35200 33562 36000 0 FreeSans 224 90 0 0 sin_out[0]
port 34 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 sin_out[1]
port 35 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 sin_outb[0]
port 36 nsew signal tristate
flabel metal2 s 9034 35200 9090 36000 0 FreeSans 224 90 0 0 sin_outb[1]
port 37 nsew signal tristate
flabel metal3 s 59200 7488 60000 7608 0 FreeSans 480 0 0 0 ud_en
port 38 nsew signal input
flabel metal4 s 8168 2128 8488 33776 0 FreeSans 1920 90 0 0 vccd1
port 39 nsew power bidirectional
flabel metal4 s 22616 2128 22936 33776 0 FreeSans 1920 90 0 0 vccd1
port 39 nsew power bidirectional
flabel metal4 s 37064 2128 37384 33776 0 FreeSans 1920 90 0 0 vccd1
port 39 nsew power bidirectional
flabel metal4 s 51512 2128 51832 33776 0 FreeSans 1920 90 0 0 vccd1
port 39 nsew power bidirectional
flabel metal4 s 15392 2128 15712 33776 0 FreeSans 1920 90 0 0 vssd1
port 40 nsew ground bidirectional
flabel metal4 s 29840 2128 30160 33776 0 FreeSans 1920 90 0 0 vssd1
port 40 nsew ground bidirectional
flabel metal4 s 44288 2128 44608 33776 0 FreeSans 1920 90 0 0 vssd1
port 40 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 36000
<< end >>
