VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO first_dual_core
  CLASS BLOCK ;
  FOREIGN first_dual_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 490.000 BY 400.000 ;
  PIN cclk_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END cclk_I[0]
  PIN cclk_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END cclk_I[1]
  PIN cclk_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 32.680 490.000 33.280 ;
    END
  END cclk_Q[0]
  PIN cclk_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 188.400 490.000 189.000 ;
    END
  END cclk_Q[1]
  PIN clk_master
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END clk_master
  PIN clk_master_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 396.000 40.850 400.000 ;
    END
  END clk_master_out
  PIN clkdiv2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END clkdiv2_I[0]
  PIN clkdiv2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END clkdiv2_I[1]
  PIN clkdiv2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 55.120 490.000 55.720 ;
    END
  END clkdiv2_Q[0]
  PIN clkdiv2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 210.840 490.000 211.440 ;
    END
  END clkdiv2_Q[1]
  PIN comp_high_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END comp_high_I[0]
  PIN comp_high_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END comp_high_I[1]
  PIN comp_high_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 77.560 490.000 78.160 ;
    END
  END comp_high_Q[0]
  PIN comp_high_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 232.600 490.000 233.200 ;
    END
  END comp_high_Q[1]
  PIN cos_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END cos_out[0]
  PIN cos_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END cos_out[1]
  PIN cos_outb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END cos_outb[0]
  PIN cos_outb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END cos_outb[1]
  PIN div2out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 396.000 95.130 400.000 ;
    END
  END div2out
  PIN fb1_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END fb1_I[0]
  PIN fb1_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END fb1_I[1]
  PIN fb1_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 121.760 490.000 122.360 ;
    END
  END fb1_Q[0]
  PIN fb1_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 277.480 490.000 278.080 ;
    END
  END fb1_Q[1]
  PIN fb2_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 396.000 476.010 400.000 ;
    END
  END fb2_I[0]
  PIN fb2_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 388.320 490.000 388.920 ;
    END
  END fb2_I[1]
  PIN fb2_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 365.880 490.000 366.480 ;
    END
  END fb2_Q[0]
  PIN fb2_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END fb2_Q[1]
  PIN gray_clk_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 396.000 367.450 400.000 ;
    END
  END gray_clk_out[10]
  PIN gray_clk_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 396.000 122.270 400.000 ;
    END
  END gray_clk_out[1]
  PIN gray_clk_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 396.000 149.410 400.000 ;
    END
  END gray_clk_out[2]
  PIN gray_clk_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 396.000 177.010 400.000 ;
    END
  END gray_clk_out[3]
  PIN gray_clk_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 396.000 204.150 400.000 ;
    END
  END gray_clk_out[4]
  PIN gray_clk_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 396.000 231.290 400.000 ;
    END
  END gray_clk_out[5]
  PIN gray_clk_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 396.000 258.430 400.000 ;
    END
  END gray_clk_out[6]
  PIN gray_clk_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 396.000 285.570 400.000 ;
    END
  END gray_clk_out[7]
  PIN gray_clk_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 396.000 312.710 400.000 ;
    END
  END gray_clk_out[8]
  PIN gray_clk_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 396.000 340.310 400.000 ;
    END
  END gray_clk_out[9]
  PIN no_ones_below_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 396.000 394.590 400.000 ;
    END
  END no_ones_below_out[0]
  PIN no_ones_below_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 396.000 421.730 400.000 ;
    END
  END no_ones_below_out[1]
  PIN no_ones_below_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 396.000 448.870 400.000 ;
    END
  END no_ones_below_out[2]
  PIN phi1b_dig_I[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END phi1b_dig_I[0]
  PIN phi1b_dig_I[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END phi1b_dig_I[1]
  PIN phi1b_dig_Q[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 99.320 490.000 99.920 ;
    END
  END phi1b_dig_Q[0]
  PIN phi1b_dig_Q[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 255.040 490.000 255.640 ;
    END
  END phi1b_dig_Q[1]
  PIN read_out_I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END read_out_I[0]
  PIN read_out_I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END read_out_I[1]
  PIN read_out_I_top[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END read_out_I_top[0]
  PIN read_out_I_top[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END read_out_I_top[1]
  PIN read_out_Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 0.000 454.850 4.000 ;
    END
  END read_out_Q[0]
  PIN read_out_Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END read_out_Q[1]
  PIN read_out_Q_top[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 321.680 490.000 322.280 ;
    END
  END read_out_Q_top[0]
  PIN read_out_Q_top[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 344.120 490.000 344.720 ;
    END
  END read_out_Q_top[1]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END rstb
  PIN rstb_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 396.000 13.710 400.000 ;
    END
  END rstb_out
  PIN sin_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 10.920 490.000 11.520 ;
    END
  END sin_out[0]
  PIN sin_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 165.960 490.000 166.560 ;
    END
  END sin_out[1]
  PIN sin_outb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 144.200 490.000 144.800 ;
    END
  END sin_outb[0]
  PIN sin_outb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 486.000 299.240 490.000 299.840 ;
    END
  END sin_outb[1]
  PIN ud_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END ud_en
  PIN ud_en_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 396.000 67.990 400.000 ;
    END
  END ud_en_out
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 389.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 484.380 389.045 ;
      LAYER met1 ;
        RECT 5.520 10.640 486.150 393.680 ;
      LAYER met2 ;
        RECT 6.990 395.720 13.150 396.965 ;
        RECT 13.990 395.720 40.290 396.965 ;
        RECT 41.130 395.720 67.430 396.965 ;
        RECT 68.270 395.720 94.570 396.965 ;
        RECT 95.410 395.720 121.710 396.965 ;
        RECT 122.550 395.720 148.850 396.965 ;
        RECT 149.690 395.720 176.450 396.965 ;
        RECT 177.290 395.720 203.590 396.965 ;
        RECT 204.430 395.720 230.730 396.965 ;
        RECT 231.570 395.720 257.870 396.965 ;
        RECT 258.710 395.720 285.010 396.965 ;
        RECT 285.850 395.720 312.150 396.965 ;
        RECT 312.990 395.720 339.750 396.965 ;
        RECT 340.590 395.720 366.890 396.965 ;
        RECT 367.730 395.720 394.030 396.965 ;
        RECT 394.870 395.720 421.170 396.965 ;
        RECT 422.010 395.720 448.310 396.965 ;
        RECT 449.150 395.720 475.450 396.965 ;
        RECT 476.290 395.720 486.120 396.965 ;
        RECT 6.990 4.280 486.120 395.720 ;
        RECT 6.990 3.670 34.770 4.280 ;
        RECT 35.610 3.670 104.690 4.280 ;
        RECT 105.530 3.670 174.610 4.280 ;
        RECT 175.450 3.670 244.530 4.280 ;
        RECT 245.370 3.670 314.450 4.280 ;
        RECT 315.290 3.670 384.370 4.280 ;
        RECT 385.210 3.670 454.290 4.280 ;
        RECT 455.130 3.670 486.120 4.280 ;
      LAYER met3 ;
        RECT 4.000 389.320 486.000 396.945 ;
        RECT 4.000 388.640 485.600 389.320 ;
        RECT 4.400 387.920 485.600 388.640 ;
        RECT 4.400 387.240 486.000 387.920 ;
        RECT 4.000 366.880 486.000 387.240 ;
        RECT 4.000 365.480 485.600 366.880 ;
        RECT 4.000 364.840 486.000 365.480 ;
        RECT 4.400 363.440 486.000 364.840 ;
        RECT 4.000 345.120 486.000 363.440 ;
        RECT 4.000 343.720 485.600 345.120 ;
        RECT 4.000 341.720 486.000 343.720 ;
        RECT 4.400 340.320 486.000 341.720 ;
        RECT 4.000 322.680 486.000 340.320 ;
        RECT 4.000 321.280 485.600 322.680 ;
        RECT 4.000 317.920 486.000 321.280 ;
        RECT 4.400 316.520 486.000 317.920 ;
        RECT 4.000 300.240 486.000 316.520 ;
        RECT 4.000 298.840 485.600 300.240 ;
        RECT 4.000 294.800 486.000 298.840 ;
        RECT 4.400 293.400 486.000 294.800 ;
        RECT 4.000 278.480 486.000 293.400 ;
        RECT 4.000 277.080 485.600 278.480 ;
        RECT 4.000 271.000 486.000 277.080 ;
        RECT 4.400 269.600 486.000 271.000 ;
        RECT 4.000 256.040 486.000 269.600 ;
        RECT 4.000 254.640 485.600 256.040 ;
        RECT 4.000 247.200 486.000 254.640 ;
        RECT 4.400 245.800 486.000 247.200 ;
        RECT 4.000 233.600 486.000 245.800 ;
        RECT 4.000 232.200 485.600 233.600 ;
        RECT 4.000 224.080 486.000 232.200 ;
        RECT 4.400 222.680 486.000 224.080 ;
        RECT 4.000 211.840 486.000 222.680 ;
        RECT 4.000 210.440 485.600 211.840 ;
        RECT 4.000 200.280 486.000 210.440 ;
        RECT 4.400 198.880 486.000 200.280 ;
        RECT 4.000 189.400 486.000 198.880 ;
        RECT 4.000 188.000 485.600 189.400 ;
        RECT 4.000 177.160 486.000 188.000 ;
        RECT 4.400 175.760 486.000 177.160 ;
        RECT 4.000 166.960 486.000 175.760 ;
        RECT 4.000 165.560 485.600 166.960 ;
        RECT 4.000 153.360 486.000 165.560 ;
        RECT 4.400 151.960 486.000 153.360 ;
        RECT 4.000 145.200 486.000 151.960 ;
        RECT 4.000 143.800 485.600 145.200 ;
        RECT 4.000 129.560 486.000 143.800 ;
        RECT 4.400 128.160 486.000 129.560 ;
        RECT 4.000 122.760 486.000 128.160 ;
        RECT 4.000 121.360 485.600 122.760 ;
        RECT 4.000 106.440 486.000 121.360 ;
        RECT 4.400 105.040 486.000 106.440 ;
        RECT 4.000 100.320 486.000 105.040 ;
        RECT 4.000 98.920 485.600 100.320 ;
        RECT 4.000 82.640 486.000 98.920 ;
        RECT 4.400 81.240 486.000 82.640 ;
        RECT 4.000 78.560 486.000 81.240 ;
        RECT 4.000 77.160 485.600 78.560 ;
        RECT 4.000 59.520 486.000 77.160 ;
        RECT 4.400 58.120 486.000 59.520 ;
        RECT 4.000 56.120 486.000 58.120 ;
        RECT 4.000 54.720 485.600 56.120 ;
        RECT 4.000 35.720 486.000 54.720 ;
        RECT 4.400 34.320 486.000 35.720 ;
        RECT 4.000 33.680 486.000 34.320 ;
        RECT 4.000 32.280 485.600 33.680 ;
        RECT 4.000 12.600 486.000 32.280 ;
        RECT 4.400 11.920 486.000 12.600 ;
        RECT 4.400 11.200 485.600 11.920 ;
        RECT 4.000 10.715 485.600 11.200 ;
      LAYER met4 ;
        RECT 68.375 389.600 469.825 396.945 ;
        RECT 68.375 66.135 97.440 389.600 ;
        RECT 99.840 66.135 174.240 389.600 ;
        RECT 176.640 66.135 251.040 389.600 ;
        RECT 253.440 66.135 327.840 389.600 ;
        RECT 330.240 66.135 404.640 389.600 ;
        RECT 407.040 66.135 469.825 389.600 ;
  END
END first_dual_core
END LIBRARY

