magic
tech sky130A
timestamp 1647840975
<< nwell >>
rect 841 -1505 3263 -1421
<< nmos >>
rect 894 -1603 909 -1561
rect 1705 -1603 1720 -1561
rect 1781 -1603 1796 -1561
rect 2575 -1603 2590 -1561
rect 2651 -1603 2666 -1561
rect 3170 -1603 3185 -1561
<< pmos >>
rect 894 -1486 909 -1444
rect 1705 -1486 1720 -1444
rect 1781 -1486 1796 -1444
rect 2575 -1486 2590 -1444
rect 2651 -1486 2666 -1444
rect 3170 -1486 3185 -1444
<< ndiff >>
rect 863 -1574 894 -1561
rect 863 -1591 869 -1574
rect 886 -1591 894 -1574
rect 863 -1603 894 -1591
rect 909 -1574 940 -1561
rect 909 -1591 916 -1574
rect 933 -1591 940 -1574
rect 909 -1603 940 -1591
rect 1674 -1574 1705 -1561
rect 1674 -1591 1680 -1574
rect 1697 -1591 1705 -1574
rect 1674 -1603 1705 -1591
rect 1720 -1573 1781 -1561
rect 1720 -1590 1745 -1573
rect 1762 -1590 1781 -1573
rect 1720 -1603 1781 -1590
rect 1796 -1574 1827 -1561
rect 1796 -1591 1803 -1574
rect 1820 -1591 1827 -1574
rect 1796 -1603 1827 -1591
rect 2544 -1574 2575 -1561
rect 2544 -1591 2550 -1574
rect 2567 -1591 2575 -1574
rect 2544 -1603 2575 -1591
rect 2590 -1573 2651 -1561
rect 2590 -1590 2615 -1573
rect 2632 -1590 2651 -1573
rect 2590 -1603 2651 -1590
rect 2666 -1574 2697 -1561
rect 2666 -1591 2673 -1574
rect 2690 -1591 2697 -1574
rect 2666 -1603 2697 -1591
rect 3139 -1574 3170 -1561
rect 3139 -1591 3145 -1574
rect 3162 -1591 3170 -1574
rect 3139 -1603 3170 -1591
rect 3185 -1574 3216 -1561
rect 3185 -1591 3192 -1574
rect 3209 -1591 3216 -1574
rect 3185 -1603 3216 -1591
<< pdiff >>
rect 863 -1456 894 -1444
rect 863 -1473 869 -1456
rect 886 -1473 894 -1456
rect 863 -1486 894 -1473
rect 909 -1456 940 -1444
rect 909 -1473 916 -1456
rect 933 -1473 940 -1456
rect 909 -1486 940 -1473
rect 1674 -1456 1705 -1444
rect 1674 -1473 1680 -1456
rect 1697 -1473 1705 -1456
rect 1674 -1486 1705 -1473
rect 1720 -1459 1781 -1444
rect 1720 -1476 1741 -1459
rect 1758 -1476 1781 -1459
rect 1720 -1486 1781 -1476
rect 1796 -1456 1827 -1444
rect 1796 -1473 1803 -1456
rect 1820 -1473 1827 -1456
rect 1796 -1486 1827 -1473
rect 2544 -1456 2575 -1444
rect 2544 -1473 2550 -1456
rect 2567 -1473 2575 -1456
rect 2544 -1486 2575 -1473
rect 2590 -1459 2651 -1444
rect 2590 -1476 2611 -1459
rect 2628 -1476 2651 -1459
rect 2590 -1486 2651 -1476
rect 2666 -1456 2697 -1444
rect 2666 -1473 2673 -1456
rect 2690 -1473 2697 -1456
rect 2666 -1486 2697 -1473
rect 3139 -1456 3170 -1444
rect 3139 -1473 3145 -1456
rect 3162 -1473 3170 -1456
rect 3139 -1486 3170 -1473
rect 3185 -1456 3216 -1444
rect 3185 -1473 3192 -1456
rect 3209 -1473 3216 -1456
rect 3185 -1486 3216 -1473
<< ndiffc >>
rect 869 -1591 886 -1574
rect 916 -1591 933 -1574
rect 1680 -1591 1697 -1574
rect 1745 -1590 1762 -1573
rect 1803 -1591 1820 -1574
rect 2550 -1591 2567 -1574
rect 2615 -1590 2632 -1573
rect 2673 -1591 2690 -1574
rect 3145 -1591 3162 -1574
rect 3192 -1591 3209 -1574
<< pdiffc >>
rect 869 -1473 886 -1456
rect 916 -1473 933 -1456
rect 1680 -1473 1697 -1456
rect 1741 -1476 1758 -1459
rect 1803 -1473 1820 -1456
rect 2550 -1473 2567 -1456
rect 2611 -1476 2628 -1459
rect 2673 -1473 2690 -1456
rect 3145 -1473 3162 -1456
rect 3192 -1473 3209 -1456
<< psubdiff >>
rect 940 -1574 969 -1561
rect 940 -1591 950 -1574
rect 967 -1591 969 -1574
rect 940 -1603 969 -1591
rect 1827 -1574 1856 -1561
rect 1827 -1591 1837 -1574
rect 1854 -1591 1856 -1574
rect 1827 -1603 1856 -1591
rect 2697 -1574 2726 -1561
rect 2697 -1591 2707 -1574
rect 2724 -1591 2726 -1574
rect 2697 -1603 2726 -1591
rect 3216 -1574 3245 -1561
rect 3216 -1591 3226 -1574
rect 3243 -1591 3245 -1574
rect 3216 -1603 3245 -1591
<< nsubdiff >>
rect 940 -1456 969 -1444
rect 940 -1473 950 -1456
rect 967 -1473 969 -1456
rect 940 -1486 969 -1473
rect 1827 -1456 1856 -1444
rect 1827 -1473 1837 -1456
rect 1854 -1473 1856 -1456
rect 1827 -1486 1856 -1473
rect 2697 -1456 2726 -1444
rect 2697 -1473 2707 -1456
rect 2724 -1473 2726 -1456
rect 2697 -1486 2726 -1473
rect 3216 -1456 3245 -1444
rect 3216 -1473 3226 -1456
rect 3243 -1473 3245 -1456
rect 3216 -1486 3245 -1473
<< psubdiffcont >>
rect 950 -1591 967 -1574
rect 1837 -1591 1854 -1574
rect 2707 -1591 2724 -1574
rect 3226 -1591 3243 -1574
<< nsubdiffcont >>
rect 950 -1473 967 -1456
rect 1837 -1473 1854 -1456
rect 2707 -1473 2724 -1456
rect 3226 -1473 3243 -1456
<< poly >>
rect 888 -1403 915 -1395
rect 1699 -1403 1726 -1395
rect 1775 -1403 1802 -1395
rect 2569 -1403 2596 -1395
rect 2645 -1403 2672 -1395
rect 3164 -1403 3191 -1395
rect 885 -1420 893 -1403
rect 910 -1420 918 -1403
rect 1696 -1420 1704 -1403
rect 1721 -1420 1729 -1403
rect 1772 -1420 1780 -1403
rect 1797 -1420 1805 -1403
rect 2566 -1420 2574 -1403
rect 2591 -1420 2599 -1403
rect 2642 -1420 2650 -1403
rect 2667 -1420 2675 -1403
rect 3161 -1420 3169 -1403
rect 3186 -1420 3194 -1403
rect 888 -1425 915 -1420
rect 1699 -1425 1726 -1420
rect 1775 -1425 1802 -1420
rect 2569 -1425 2596 -1420
rect 2645 -1425 2672 -1420
rect 3164 -1425 3191 -1420
rect 894 -1444 909 -1425
rect 1705 -1444 1720 -1425
rect 1781 -1444 1796 -1425
rect 2575 -1444 2590 -1425
rect 2651 -1444 2666 -1425
rect 3170 -1444 3185 -1425
rect 894 -1499 909 -1486
rect 1705 -1499 1720 -1486
rect 1781 -1499 1796 -1486
rect 2575 -1499 2590 -1486
rect 2651 -1499 2666 -1486
rect 3170 -1499 3185 -1486
rect 894 -1561 909 -1548
rect 1705 -1561 1720 -1548
rect 1781 -1561 1796 -1548
rect 2575 -1561 2590 -1548
rect 2651 -1561 2666 -1548
rect 3170 -1561 3185 -1548
rect 894 -1619 909 -1603
rect 1705 -1619 1720 -1603
rect 1781 -1619 1796 -1603
rect 2575 -1619 2590 -1603
rect 2651 -1619 2666 -1603
rect 3170 -1619 3185 -1603
rect 888 -1624 915 -1619
rect 1699 -1624 1726 -1619
rect 1775 -1624 1802 -1619
rect 2569 -1624 2596 -1619
rect 2645 -1624 2672 -1619
rect 3164 -1624 3191 -1619
rect 885 -1641 893 -1624
rect 910 -1641 918 -1624
rect 1696 -1641 1704 -1624
rect 1721 -1641 1729 -1624
rect 1772 -1641 1780 -1624
rect 1797 -1641 1805 -1624
rect 2566 -1641 2574 -1624
rect 2591 -1641 2599 -1624
rect 2642 -1641 2650 -1624
rect 2667 -1641 2675 -1624
rect 3161 -1641 3169 -1624
rect 3186 -1641 3194 -1624
rect 888 -1649 915 -1641
rect 1699 -1649 1726 -1641
rect 1775 -1649 1802 -1641
rect 2569 -1649 2596 -1641
rect 2645 -1649 2672 -1641
rect 3164 -1649 3191 -1641
<< polycont >>
rect 893 -1420 910 -1403
rect 1704 -1420 1721 -1403
rect 1780 -1420 1797 -1403
rect 2574 -1420 2591 -1403
rect 2650 -1420 2667 -1403
rect 3169 -1420 3186 -1403
rect 893 -1641 910 -1624
rect 1704 -1641 1721 -1624
rect 1780 -1641 1797 -1624
rect 2574 -1641 2591 -1624
rect 2650 -1641 2667 -1624
rect 3169 -1641 3186 -1624
<< locali >>
rect 944 -1367 950 -1350
rect 967 -1367 972 -1350
rect 885 -1420 893 -1403
rect 910 -1420 918 -1403
rect 869 -1456 886 -1448
rect 869 -1517 886 -1473
rect 869 -1574 886 -1534
rect 869 -1599 886 -1591
rect 916 -1456 933 -1448
rect 916 -1520 933 -1473
rect 950 -1456 967 -1367
rect 1704 -1403 1721 -1287
rect 1780 -1308 1797 -1304
rect 1780 -1403 1797 -1325
rect 1837 -1350 1854 -1347
rect 1834 -1367 1837 -1350
rect 1854 -1367 1857 -1350
rect 1696 -1420 1704 -1403
rect 1721 -1420 1729 -1403
rect 1772 -1420 1780 -1403
rect 1797 -1420 1805 -1403
rect 950 -1481 967 -1473
rect 1680 -1456 1697 -1448
rect 1680 -1517 1697 -1473
rect 916 -1537 924 -1520
rect 916 -1574 933 -1537
rect 916 -1599 933 -1591
rect 950 -1574 967 -1566
rect 893 -1624 910 -1621
rect 885 -1641 893 -1624
rect 910 -1641 918 -1624
rect 893 -1644 910 -1641
rect 950 -1683 967 -1591
rect 1680 -1574 1697 -1534
rect 1680 -1599 1697 -1591
rect 1727 -1459 1773 -1448
rect 1727 -1476 1741 -1459
rect 1758 -1476 1773 -1459
rect 1727 -1521 1773 -1476
rect 1744 -1538 1773 -1521
rect 1727 -1573 1773 -1538
rect 1727 -1590 1745 -1573
rect 1762 -1590 1773 -1573
rect 1727 -1599 1773 -1590
rect 1803 -1456 1820 -1448
rect 1803 -1520 1820 -1473
rect 1837 -1456 1854 -1367
rect 2574 -1403 2591 -1287
rect 2650 -1403 2667 -1321
rect 2707 -1350 2724 -1347
rect 2704 -1367 2707 -1350
rect 2724 -1367 2727 -1350
rect 2566 -1420 2574 -1403
rect 2591 -1420 2599 -1403
rect 2642 -1420 2650 -1403
rect 2667 -1420 2675 -1403
rect 1837 -1481 1854 -1473
rect 2550 -1456 2567 -1448
rect 2550 -1517 2567 -1473
rect 1803 -1537 1811 -1520
rect 1803 -1574 1820 -1537
rect 1803 -1599 1820 -1591
rect 1837 -1574 1854 -1566
rect 1696 -1641 1704 -1624
rect 1721 -1641 1729 -1624
rect 1772 -1641 1780 -1624
rect 1797 -1641 1805 -1624
rect 1704 -1765 1721 -1641
rect 1780 -1722 1797 -1641
rect 1837 -1683 1854 -1591
rect 2550 -1574 2567 -1534
rect 2550 -1599 2567 -1591
rect 2597 -1459 2643 -1448
rect 2597 -1476 2611 -1459
rect 2628 -1476 2643 -1459
rect 2597 -1521 2643 -1476
rect 2614 -1538 2643 -1521
rect 2597 -1573 2643 -1538
rect 2597 -1590 2615 -1573
rect 2632 -1590 2643 -1573
rect 2597 -1599 2643 -1590
rect 2673 -1456 2690 -1448
rect 2673 -1520 2690 -1473
rect 2707 -1456 2724 -1367
rect 3169 -1403 3186 -1287
rect 3226 -1350 3243 -1347
rect 3223 -1367 3226 -1350
rect 3243 -1367 3246 -1350
rect 3161 -1420 3169 -1403
rect 3186 -1420 3194 -1403
rect 2707 -1481 2724 -1473
rect 3145 -1456 3162 -1448
rect 3145 -1519 3162 -1473
rect 2673 -1537 2681 -1520
rect 3153 -1536 3162 -1519
rect 2673 -1574 2690 -1537
rect 2673 -1599 2690 -1591
rect 2707 -1574 2724 -1566
rect 2566 -1641 2574 -1624
rect 2591 -1641 2599 -1624
rect 2642 -1641 2650 -1624
rect 2667 -1641 2675 -1624
rect 1780 -1748 1797 -1739
rect 2574 -1765 2591 -1641
rect 2650 -1731 2667 -1641
rect 2707 -1683 2724 -1591
rect 3145 -1574 3162 -1536
rect 3145 -1599 3162 -1591
rect 3192 -1456 3209 -1448
rect 3192 -1520 3209 -1473
rect 3226 -1456 3243 -1367
rect 3226 -1481 3243 -1473
rect 3192 -1537 3200 -1520
rect 3192 -1574 3209 -1537
rect 3192 -1599 3209 -1591
rect 3226 -1574 3243 -1566
rect 3161 -1641 3169 -1624
rect 3186 -1641 3194 -1624
rect 2724 -1700 2730 -1683
rect 3169 -1765 3186 -1641
rect 3226 -1683 3243 -1591
<< viali >>
rect 1704 -1287 1721 -1270
rect 950 -1367 967 -1350
rect 893 -1420 910 -1403
rect 869 -1534 886 -1517
rect 2574 -1287 2591 -1270
rect 1780 -1325 1797 -1308
rect 1837 -1367 1854 -1350
rect 924 -1537 941 -1520
rect 1680 -1534 1697 -1517
rect 893 -1641 910 -1624
rect 1727 -1538 1744 -1521
rect 3169 -1287 3186 -1270
rect 2650 -1321 2667 -1304
rect 2707 -1367 2724 -1350
rect 1811 -1537 1828 -1520
rect 2550 -1534 2567 -1517
rect 950 -1700 967 -1683
rect 2597 -1538 2614 -1521
rect 3226 -1367 3243 -1350
rect 2681 -1537 2698 -1520
rect 3136 -1536 3153 -1519
rect 1837 -1700 1854 -1683
rect 1780 -1739 1797 -1722
rect 1704 -1782 1721 -1765
rect 3200 -1537 3217 -1520
rect 2707 -1700 2724 -1683
rect 2650 -1748 2667 -1731
rect 2574 -1782 2591 -1765
rect 3226 -1700 3243 -1683
rect 3169 -1782 3186 -1765
<< metal1 >>
rect 1698 -1270 1727 -1264
rect 1698 -1287 1704 -1270
rect 1721 -1273 1727 -1270
rect 2568 -1270 2597 -1264
rect 2568 -1273 2574 -1270
rect 1721 -1287 2574 -1273
rect 2591 -1273 2597 -1270
rect 3163 -1270 3192 -1267
rect 3163 -1273 3169 -1270
rect 2591 -1287 3169 -1273
rect 3186 -1273 3192 -1270
rect 3186 -1287 5596 -1273
rect 1698 -1290 1727 -1287
rect 2568 -1290 2597 -1287
rect 3163 -1290 3192 -1287
rect 2644 -1304 2672 -1301
rect 893 -1308 2650 -1304
rect 893 -1318 1780 -1308
rect 893 -1397 910 -1318
rect 1774 -1325 1780 -1318
rect 1797 -1318 2650 -1308
rect 1797 -1325 1803 -1318
rect 1774 -1330 1803 -1325
rect 2644 -1321 2650 -1318
rect 2667 -1318 5596 -1304
rect 2667 -1321 2672 -1318
rect 2644 -1327 2672 -1321
rect 947 -1350 970 -1347
rect 1834 -1350 1857 -1347
rect 2704 -1350 2727 -1347
rect 3223 -1350 3246 -1347
rect 944 -1367 950 -1350
rect 967 -1367 1837 -1350
rect 1854 -1367 2707 -1350
rect 2724 -1367 3226 -1350
rect 3243 -1367 5596 -1350
rect 947 -1370 970 -1367
rect 1834 -1370 1857 -1367
rect 2704 -1370 2727 -1367
rect 3223 -1370 3246 -1367
rect 889 -1403 914 -1397
rect 889 -1420 893 -1403
rect 910 -1420 914 -1403
rect 889 -1426 914 -1420
rect 862 -1512 892 -1511
rect 859 -1514 902 -1512
rect 859 -1540 864 -1514
rect 890 -1540 902 -1514
rect 978 -1516 1008 -1515
rect 916 -1518 1011 -1516
rect 916 -1520 980 -1518
rect 916 -1537 924 -1520
rect 941 -1537 980 -1520
rect 916 -1540 980 -1537
rect 859 -1549 902 -1540
rect 968 -1544 980 -1540
rect 1006 -1544 1011 -1518
rect 968 -1553 1011 -1544
rect 1633 -1517 1700 -1509
rect 1722 -1516 1756 -1513
rect 1865 -1516 1895 -1515
rect 1633 -1518 1680 -1517
rect 1633 -1544 1638 -1518
rect 1664 -1534 1680 -1518
rect 1697 -1534 1700 -1517
rect 1664 -1544 1700 -1534
rect 1633 -1546 1700 -1544
rect 1721 -1518 1756 -1516
rect 1721 -1544 1724 -1518
rect 1750 -1544 1756 -1518
rect 1803 -1518 1898 -1516
rect 1803 -1520 1867 -1518
rect 1803 -1537 1811 -1520
rect 1828 -1537 1867 -1520
rect 1803 -1540 1867 -1537
rect 1721 -1546 1756 -1544
rect 1636 -1547 1666 -1546
rect 1722 -1549 1756 -1546
rect 1855 -1544 1867 -1540
rect 1893 -1544 1898 -1518
rect 1855 -1553 1898 -1544
rect 2503 -1517 2570 -1509
rect 2592 -1516 2626 -1513
rect 2735 -1516 2765 -1515
rect 2503 -1518 2550 -1517
rect 2503 -1544 2508 -1518
rect 2534 -1534 2550 -1518
rect 2567 -1534 2570 -1517
rect 2534 -1544 2570 -1534
rect 2503 -1546 2570 -1544
rect 2591 -1518 2626 -1516
rect 2591 -1544 2594 -1518
rect 2620 -1544 2626 -1518
rect 2673 -1518 2768 -1516
rect 2673 -1520 2737 -1518
rect 2673 -1537 2681 -1520
rect 2698 -1537 2737 -1520
rect 2673 -1540 2737 -1537
rect 2591 -1546 2626 -1544
rect 2506 -1547 2536 -1546
rect 2592 -1549 2626 -1546
rect 2725 -1544 2737 -1540
rect 2763 -1544 2768 -1518
rect 2725 -1553 2768 -1544
rect 3120 -1518 3163 -1509
rect 3254 -1516 3284 -1515
rect 3120 -1544 3125 -1518
rect 3151 -1519 3163 -1518
rect 3153 -1536 3163 -1519
rect 3151 -1544 3163 -1536
rect 3192 -1518 3287 -1516
rect 3192 -1520 3256 -1518
rect 3192 -1537 3200 -1520
rect 3217 -1537 3256 -1520
rect 3192 -1540 3256 -1537
rect 3120 -1546 3163 -1544
rect 3244 -1544 3256 -1540
rect 3282 -1544 3287 -1518
rect 3123 -1547 3153 -1546
rect 3244 -1553 3287 -1544
rect 5496 -1579 5523 -1576
rect 5523 -1599 5596 -1585
rect 5496 -1608 5523 -1605
rect 890 -1624 913 -1618
rect 890 -1641 893 -1624
rect 910 -1641 913 -1624
rect 890 -1644 913 -1641
rect 893 -1734 910 -1644
rect 945 -1677 972 -1675
rect 1832 -1677 1859 -1675
rect 2702 -1677 2729 -1675
rect 3221 -1677 3248 -1675
rect 944 -1678 973 -1677
rect 944 -1705 945 -1678
rect 972 -1705 973 -1678
rect 944 -1706 973 -1705
rect 1831 -1678 1860 -1677
rect 1831 -1705 1832 -1678
rect 1859 -1705 1860 -1678
rect 1831 -1706 1860 -1705
rect 2701 -1678 2730 -1677
rect 2701 -1705 2702 -1678
rect 2729 -1705 2730 -1678
rect 2701 -1706 2730 -1705
rect 3220 -1678 3249 -1677
rect 3220 -1705 3221 -1678
rect 3248 -1705 3249 -1678
rect 3220 -1706 3249 -1705
rect 945 -1708 972 -1706
rect 1832 -1708 1859 -1706
rect 2702 -1708 2729 -1706
rect 3221 -1708 3248 -1706
rect 1771 -1722 1803 -1714
rect 1771 -1734 1780 -1722
rect 893 -1739 1780 -1734
rect 1797 -1734 1803 -1722
rect 2644 -1731 2673 -1724
rect 2644 -1734 2650 -1731
rect 1797 -1739 2650 -1734
rect 893 -1748 2650 -1739
rect 2667 -1734 2673 -1731
rect 2667 -1748 5596 -1734
rect 2644 -1752 2673 -1748
rect 1698 -1765 1727 -1762
rect 1698 -1782 1704 -1765
rect 1721 -1766 1727 -1765
rect 2568 -1765 2598 -1762
rect 2568 -1766 2574 -1765
rect 1721 -1780 2574 -1766
rect 1721 -1782 1727 -1780
rect 1698 -1788 1727 -1782
rect 2568 -1782 2574 -1780
rect 2591 -1766 2598 -1765
rect 3163 -1765 3192 -1762
rect 3163 -1766 3169 -1765
rect 2591 -1780 3169 -1766
rect 2591 -1782 2598 -1780
rect 2568 -1791 2598 -1782
rect 3163 -1782 3169 -1780
rect 3186 -1766 3192 -1765
rect 3186 -1780 5596 -1766
rect 3186 -1782 3192 -1780
rect 3163 -1788 3192 -1782
<< via1 >>
rect 864 -1517 890 -1514
rect 864 -1534 869 -1517
rect 869 -1534 886 -1517
rect 886 -1534 890 -1517
rect 864 -1540 890 -1534
rect 980 -1544 1006 -1518
rect 1638 -1544 1664 -1518
rect 1724 -1521 1750 -1518
rect 1724 -1538 1727 -1521
rect 1727 -1538 1744 -1521
rect 1744 -1538 1750 -1521
rect 1724 -1544 1750 -1538
rect 1867 -1544 1893 -1518
rect 2508 -1544 2534 -1518
rect 2594 -1521 2620 -1518
rect 2594 -1538 2597 -1521
rect 2597 -1538 2614 -1521
rect 2614 -1538 2620 -1521
rect 2594 -1544 2620 -1538
rect 2737 -1544 2763 -1518
rect 3125 -1519 3151 -1518
rect 3125 -1536 3136 -1519
rect 3136 -1536 3151 -1519
rect 3125 -1544 3151 -1536
rect 3256 -1544 3282 -1518
rect 5496 -1605 5523 -1579
rect 945 -1683 972 -1678
rect 945 -1700 950 -1683
rect 950 -1700 967 -1683
rect 967 -1700 972 -1683
rect 945 -1705 972 -1700
rect 1832 -1683 1859 -1678
rect 1832 -1700 1837 -1683
rect 1837 -1700 1854 -1683
rect 1854 -1700 1859 -1683
rect 1832 -1705 1859 -1700
rect 2702 -1683 2729 -1678
rect 2702 -1700 2707 -1683
rect 2707 -1700 2724 -1683
rect 2724 -1700 2729 -1683
rect 2702 -1705 2729 -1700
rect 3221 -1683 3248 -1678
rect 3221 -1700 3226 -1683
rect 3226 -1700 3243 -1683
rect 3243 -1700 3248 -1683
rect 3221 -1705 3248 -1700
<< metal2 >>
rect 859 -1513 895 -1508
rect 859 -1541 863 -1513
rect 891 -1541 895 -1513
rect 859 -1546 895 -1541
rect 975 -1517 1011 -1512
rect 975 -1545 979 -1517
rect 1007 -1545 1011 -1517
rect 975 -1550 1011 -1545
rect 1633 -1517 1669 -1512
rect 1633 -1545 1637 -1517
rect 1665 -1545 1669 -1517
rect 1633 -1550 1669 -1545
rect 1718 -1517 1756 -1513
rect 1718 -1545 1723 -1517
rect 1751 -1545 1756 -1517
rect 1718 -1549 1756 -1545
rect 1862 -1517 1898 -1512
rect 1862 -1545 1866 -1517
rect 1894 -1545 1898 -1517
rect 1862 -1550 1898 -1545
rect 2503 -1517 2539 -1512
rect 2503 -1545 2507 -1517
rect 2535 -1545 2539 -1517
rect 2503 -1550 2539 -1545
rect 2588 -1517 2626 -1513
rect 2588 -1545 2593 -1517
rect 2621 -1545 2626 -1517
rect 2588 -1549 2626 -1545
rect 2732 -1517 2768 -1512
rect 2732 -1545 2736 -1517
rect 2764 -1545 2768 -1517
rect 2732 -1550 2768 -1545
rect 3120 -1517 3156 -1512
rect 3120 -1545 3124 -1517
rect 3152 -1545 3156 -1517
rect 3120 -1550 3156 -1545
rect 3251 -1517 3287 -1512
rect 3251 -1545 3255 -1517
rect 3283 -1545 3287 -1517
rect 3251 -1550 3287 -1545
rect 5492 -1575 5526 -1570
rect 5492 -1614 5526 -1609
rect 945 -1678 972 -1675
rect 1832 -1678 1859 -1675
rect 2702 -1678 2729 -1675
rect 3221 -1678 3248 -1675
rect 940 -1706 945 -1678
rect 973 -1706 978 -1678
rect 1827 -1706 1832 -1678
rect 1860 -1706 1865 -1678
rect 2697 -1706 2702 -1678
rect 2730 -1706 2735 -1678
rect 3216 -1706 3221 -1678
rect 3249 -1706 3254 -1678
rect 945 -1708 972 -1706
rect 1832 -1708 1859 -1706
rect 2702 -1708 2729 -1706
rect 3221 -1708 3248 -1706
<< via2 >>
rect 863 -1514 891 -1513
rect 863 -1540 864 -1514
rect 864 -1540 890 -1514
rect 890 -1540 891 -1514
rect 863 -1541 891 -1540
rect 979 -1518 1007 -1517
rect 979 -1544 980 -1518
rect 980 -1544 1006 -1518
rect 1006 -1544 1007 -1518
rect 979 -1545 1007 -1544
rect 1637 -1518 1665 -1517
rect 1637 -1544 1638 -1518
rect 1638 -1544 1664 -1518
rect 1664 -1544 1665 -1518
rect 1637 -1545 1665 -1544
rect 1723 -1518 1751 -1517
rect 1723 -1544 1724 -1518
rect 1724 -1544 1750 -1518
rect 1750 -1544 1751 -1518
rect 1723 -1545 1751 -1544
rect 1866 -1518 1894 -1517
rect 1866 -1544 1867 -1518
rect 1867 -1544 1893 -1518
rect 1893 -1544 1894 -1518
rect 1866 -1545 1894 -1544
rect 2507 -1518 2535 -1517
rect 2507 -1544 2508 -1518
rect 2508 -1544 2534 -1518
rect 2534 -1544 2535 -1518
rect 2507 -1545 2535 -1544
rect 2593 -1518 2621 -1517
rect 2593 -1544 2594 -1518
rect 2594 -1544 2620 -1518
rect 2620 -1544 2621 -1518
rect 2593 -1545 2621 -1544
rect 2736 -1518 2764 -1517
rect 2736 -1544 2737 -1518
rect 2737 -1544 2763 -1518
rect 2763 -1544 2764 -1518
rect 2736 -1545 2764 -1544
rect 3124 -1518 3152 -1517
rect 3124 -1544 3125 -1518
rect 3125 -1544 3151 -1518
rect 3151 -1544 3152 -1518
rect 3124 -1545 3152 -1544
rect 3255 -1518 3283 -1517
rect 3255 -1544 3256 -1518
rect 3256 -1544 3282 -1518
rect 3282 -1544 3283 -1518
rect 3255 -1545 3283 -1544
rect 5492 -1579 5526 -1575
rect 5492 -1605 5496 -1579
rect 5496 -1605 5523 -1579
rect 5523 -1605 5526 -1579
rect 5492 -1609 5526 -1605
rect 945 -1705 972 -1678
rect 972 -1705 973 -1678
rect 945 -1706 973 -1705
rect 1832 -1705 1859 -1678
rect 1859 -1705 1860 -1678
rect 1832 -1706 1860 -1705
rect 2702 -1705 2729 -1678
rect 2729 -1705 2730 -1678
rect 2702 -1706 2730 -1705
rect 3221 -1705 3248 -1678
rect 3248 -1705 3249 -1678
rect 3221 -1706 3249 -1705
<< metal3 >>
rect -2644 2790 -2315 2853
rect -2644 2758 -2580 2790
rect -2548 2758 -2315 2790
rect -2644 2690 -2315 2758
rect -2483 2627 -2172 2690
rect -2483 2595 -2252 2627
rect -2220 2595 -2172 2627
rect -2483 2527 -2172 2595
rect -2644 2464 -2315 2527
rect -2644 2432 -2580 2464
rect -2548 2432 -2315 2464
rect -2644 2364 -2315 2432
rect -2483 2301 -2172 2364
rect -2483 2269 -2252 2301
rect -2220 2269 -2172 2301
rect -2483 2201 -2172 2269
rect -2644 2138 -2315 2201
rect -2644 2106 -2580 2138
rect -2548 2106 -2315 2138
rect -2644 2038 -2315 2106
rect -2483 1975 -2172 2038
rect -2483 1943 -2252 1975
rect -2220 1943 -2172 1975
rect -2483 1875 -2172 1943
rect -2644 1812 -2315 1875
rect -2644 1780 -2580 1812
rect -2548 1780 -2315 1812
rect -2644 1712 -2315 1780
rect -2483 1649 -2172 1712
rect -2483 1617 -2252 1649
rect -2220 1617 -2172 1649
rect -2483 1549 -2172 1617
rect -2644 1486 -2315 1549
rect -2644 1454 -2580 1486
rect -2548 1454 -2315 1486
rect -2644 1386 -2315 1454
rect -2483 1323 -2172 1386
rect -2483 1291 -2252 1323
rect -2220 1291 -2172 1323
rect -2483 1223 -2172 1291
rect -2644 1160 -2315 1223
rect -2644 1128 -2580 1160
rect -2548 1128 -2315 1160
rect -2644 1060 -2315 1128
rect -2483 997 -2172 1060
rect -2483 965 -2252 997
rect -2220 965 -2172 997
rect -2483 897 -2172 965
rect -2644 834 -2315 897
rect -2644 802 -2580 834
rect -2548 802 -2315 834
rect -2644 734 -2315 802
rect -2483 671 -2172 734
rect -2483 639 -2252 671
rect -2220 639 -2172 671
rect -2483 571 -2172 639
rect -2644 508 -2315 571
rect -2644 476 -2580 508
rect -2548 476 -2315 508
rect -2644 408 -2315 476
rect -2483 345 -2172 408
rect -2483 313 -2252 345
rect -2220 313 -2172 345
rect -2483 245 -2172 313
rect -2644 182 -2315 245
rect -2644 150 -2580 182
rect -2548 150 -2315 182
rect -2644 82 -2315 150
rect -2483 19 -2172 82
rect -2483 -13 -2252 19
rect -2220 -13 -2172 19
rect -2483 -81 -2172 -13
rect -2644 -144 -2315 -81
rect -2644 -176 -2580 -144
rect -2548 -176 -2315 -144
rect -2644 -244 -2315 -176
rect -2483 -307 -2172 -244
rect -2483 -339 -2252 -307
rect -2220 -339 -2172 -307
rect -2483 -407 -2172 -339
rect -2644 -470 -2315 -407
rect -2644 -502 -2580 -470
rect -2548 -502 -2315 -470
rect -2644 -570 -2315 -502
rect -2483 -633 -2172 -570
rect -2483 -665 -2252 -633
rect -2220 -665 -2172 -633
rect -2483 -733 -2172 -665
rect -2644 -796 -2315 -733
rect -2644 -828 -2580 -796
rect -2548 -828 -2315 -796
rect -2644 -896 -2315 -828
rect -2483 -897 -2315 -896
rect -2483 -960 -2172 -897
rect -2483 -992 -2252 -960
rect -2220 -992 -2172 -960
rect -2483 -1060 -2172 -992
rect -2644 -1123 -2315 -1060
rect -2644 -1155 -2580 -1123
rect -2548 -1155 -2315 -1123
rect -2644 -1223 -2315 -1155
rect -2483 -1387 -2315 -1223
rect -2092 -1250 5604 2862
rect -2644 -1443 -2315 -1387
rect 1057 -1306 1149 -1250
rect -2644 -1450 782 -1443
rect -2644 -1482 -2580 -1450
rect -2548 -1482 782 -1450
rect -2644 -1550 782 -1482
rect 853 -1511 902 -1501
rect 853 -1543 861 -1511
rect 893 -1543 902 -1511
rect 853 -1549 902 -1543
rect -2483 -1579 782 -1550
rect 858 -1553 902 -1549
rect 968 -1515 1017 -1505
rect 968 -1547 977 -1515
rect 1009 -1547 1017 -1515
rect 968 -1557 1017 -1547
rect -2483 -1583 828 -1579
rect -2483 -1609 839 -1583
rect 798 -1667 839 -1609
rect 1057 -1667 1585 -1306
rect 1627 -1515 1676 -1505
rect 1627 -1547 1635 -1515
rect 1667 -1547 1676 -1515
rect 1627 -1557 1676 -1547
rect 1711 -1515 1763 -1507
rect 1711 -1547 1721 -1515
rect 1753 -1547 1763 -1515
rect 1711 -1556 1763 -1547
rect 1855 -1515 1904 -1505
rect 1855 -1547 1864 -1515
rect 1896 -1547 1904 -1515
rect 1855 -1557 1904 -1547
rect 1936 -1667 2464 -1430
rect 2497 -1515 2546 -1505
rect 2497 -1547 2505 -1515
rect 2537 -1547 2546 -1515
rect 2497 -1557 2546 -1547
rect 2581 -1515 2633 -1507
rect 2581 -1547 2591 -1515
rect 2623 -1547 2633 -1515
rect 2581 -1556 2633 -1547
rect 2725 -1515 2774 -1505
rect 2725 -1547 2734 -1515
rect 2766 -1547 2774 -1515
rect 2725 -1557 2774 -1547
rect 2806 -1667 3084 -1423
rect 3114 -1515 3163 -1505
rect 3114 -1547 3122 -1515
rect 3154 -1547 3163 -1515
rect 3114 -1557 3163 -1547
rect 3244 -1515 3293 -1505
rect 3244 -1547 3253 -1515
rect 3285 -1547 3293 -1515
rect 3244 -1551 3293 -1547
rect 3244 -1557 3286 -1551
rect 5428 -1575 5592 -1502
rect 5428 -1609 5492 -1575
rect 5526 -1609 5592 -1575
rect 798 -1678 3255 -1667
rect 798 -1706 945 -1678
rect 973 -1706 1832 -1678
rect 1860 -1706 2702 -1678
rect 2730 -1706 3221 -1678
rect 3249 -1706 3255 -1678
rect 798 -1716 3255 -1706
rect 1057 -1734 1585 -1716
rect 1057 -1797 1151 -1734
rect 5428 -1797 5592 -1609
rect -2093 -4825 3019 -1797
rect 3075 -4825 5604 -1797
<< via3 >>
rect -2580 2758 -2548 2790
rect -2252 2595 -2220 2627
rect -2580 2432 -2548 2464
rect -2252 2269 -2220 2301
rect -2580 2106 -2548 2138
rect -2252 1943 -2220 1975
rect -2580 1780 -2548 1812
rect -2252 1617 -2220 1649
rect -2580 1454 -2548 1486
rect -2252 1291 -2220 1323
rect -2580 1128 -2548 1160
rect -2252 965 -2220 997
rect -2580 802 -2548 834
rect -2252 639 -2220 671
rect -2580 476 -2548 508
rect -2252 313 -2220 345
rect -2580 150 -2548 182
rect -2252 -13 -2220 19
rect -2580 -176 -2548 -144
rect -2252 -339 -2220 -307
rect -2580 -502 -2548 -470
rect -2252 -665 -2220 -633
rect -2580 -828 -2548 -796
rect -2252 -992 -2220 -960
rect -2580 -1155 -2548 -1123
rect -2580 -1482 -2548 -1450
rect 861 -1513 893 -1511
rect 861 -1541 863 -1513
rect 863 -1541 891 -1513
rect 891 -1541 893 -1513
rect 861 -1543 893 -1541
rect 977 -1517 1009 -1515
rect 977 -1545 979 -1517
rect 979 -1545 1007 -1517
rect 1007 -1545 1009 -1517
rect 977 -1547 1009 -1545
rect 1635 -1517 1667 -1515
rect 1635 -1545 1637 -1517
rect 1637 -1545 1665 -1517
rect 1665 -1545 1667 -1517
rect 1635 -1547 1667 -1545
rect 1721 -1517 1753 -1515
rect 1721 -1545 1723 -1517
rect 1723 -1545 1751 -1517
rect 1751 -1545 1753 -1517
rect 1721 -1547 1753 -1545
rect 1864 -1517 1896 -1515
rect 1864 -1545 1866 -1517
rect 1866 -1545 1894 -1517
rect 1894 -1545 1896 -1517
rect 1864 -1547 1896 -1545
rect 2505 -1517 2537 -1515
rect 2505 -1545 2507 -1517
rect 2507 -1545 2535 -1517
rect 2535 -1545 2537 -1517
rect 2505 -1547 2537 -1545
rect 2591 -1517 2623 -1515
rect 2591 -1545 2593 -1517
rect 2593 -1545 2621 -1517
rect 2621 -1545 2623 -1517
rect 2591 -1547 2623 -1545
rect 2734 -1517 2766 -1515
rect 2734 -1545 2736 -1517
rect 2736 -1545 2764 -1517
rect 2764 -1545 2766 -1517
rect 2734 -1547 2766 -1545
rect 3122 -1517 3154 -1515
rect 3122 -1545 3124 -1517
rect 3124 -1545 3152 -1517
rect 3152 -1545 3154 -1517
rect 3122 -1547 3154 -1545
rect 3253 -1517 3285 -1515
rect 3253 -1545 3255 -1517
rect 3255 -1545 3283 -1517
rect 3283 -1545 3285 -1517
rect 3253 -1547 3285 -1545
rect 5492 -1609 5526 -1575
<< mimcap >>
rect -2078 1187 922 2848
rect -2078 1069 757 1187
rect 875 1069 922 1187
rect -2078 848 922 1069
rect 1006 1184 4006 2848
rect 1006 1066 1059 1184
rect 1177 1161 4006 1184
rect 1177 1066 3847 1161
rect 1006 1043 3847 1066
rect 3965 1043 4006 1161
rect 1006 848 4006 1043
rect 4090 1194 5590 2848
rect 4090 1076 4143 1194
rect 4261 1076 5590 1194
rect 4090 848 5590 1076
rect -2078 540 922 764
rect -2078 422 767 540
rect 885 422 922 540
rect -2078 -1071 922 422
rect -2078 -1189 -1858 -1071
rect -1740 -1189 922 -1071
rect -2078 -1236 922 -1189
rect 1006 547 4006 764
rect 1006 429 1040 547
rect 1158 505 4006 547
rect 1158 429 3825 505
rect 1006 387 3825 429
rect 3943 387 4006 505
rect 1006 -1236 4006 387
rect 4090 488 5590 764
rect 4090 370 4133 488
rect 4251 370 5590 488
rect 4090 -1236 5590 370
rect 1071 -1514 1571 -1320
rect 1071 -1549 1091 -1514
rect 1127 -1549 1519 -1514
rect 1071 -1550 1519 -1549
rect 1553 -1550 1571 -1514
rect 1071 -1720 1571 -1550
rect 1950 -1512 2450 -1444
rect 1950 -1548 1965 -1512
rect 2000 -1515 2450 -1512
rect 2000 -1548 2405 -1515
rect 1950 -1549 2405 -1548
rect 2440 -1549 2450 -1515
rect 1950 -1644 2450 -1549
rect 2820 -1513 3070 -1437
rect 2820 -1547 2830 -1513
rect 2864 -1515 3070 -1513
rect 2864 -1547 3026 -1515
rect 2820 -1550 3026 -1547
rect 3060 -1550 3070 -1515
rect 2820 -1637 3070 -1550
rect -2079 -1864 421 -1811
rect -2079 -1982 -1843 -1864
rect -1725 -1982 421 -1864
rect -2079 -4811 421 -1982
rect 505 -1847 3005 -1811
rect 505 -1965 725 -1847
rect 843 -1965 3005 -1847
rect 505 -4811 3005 -1965
rect 3089 -1864 5590 -1811
rect 3089 -1982 3327 -1864
rect 3445 -1982 5590 -1864
rect 3089 -4811 5590 -1982
<< mimcapcontact >>
rect 757 1069 875 1187
rect 1059 1066 1177 1184
rect 3847 1043 3965 1161
rect 4143 1076 4261 1194
rect 767 422 885 540
rect -1858 -1189 -1740 -1071
rect 1040 429 1158 547
rect 3825 387 3943 505
rect 4133 370 4251 488
rect 1091 -1549 1127 -1514
rect 1519 -1550 1553 -1514
rect 1965 -1548 2000 -1512
rect 2405 -1549 2440 -1515
rect 2830 -1547 2864 -1513
rect 3026 -1550 3060 -1515
rect -1843 -1982 -1725 -1864
rect 725 -1965 843 -1847
rect 3327 -1982 3445 -1864
<< metal4 >>
rect -2644 2834 -2493 2853
rect -2644 2716 -2622 2834
rect -2504 2716 -2493 2834
rect -2644 2690 -2493 2716
rect -2644 2508 -2493 2527
rect -2644 2390 -2622 2508
rect -2504 2390 -2493 2508
rect -2644 2364 -2493 2390
rect -2644 2182 -2493 2201
rect -2644 2064 -2622 2182
rect -2504 2064 -2493 2182
rect -2644 2038 -2493 2064
rect -2644 1856 -2493 1875
rect -2644 1738 -2622 1856
rect -2504 1738 -2493 1856
rect -2644 1712 -2493 1738
rect -2644 1530 -2493 1549
rect -2644 1412 -2622 1530
rect -2504 1412 -2493 1530
rect -2644 1386 -2493 1412
rect -2644 1204 -2493 1223
rect -2644 1086 -2622 1204
rect -2504 1086 -2493 1204
rect -2644 1060 -2493 1086
rect -2644 878 -2493 897
rect -2644 760 -2622 878
rect -2504 760 -2493 878
rect -2644 734 -2493 760
rect -2644 552 -2493 571
rect -2644 434 -2622 552
rect -2504 434 -2493 552
rect -2644 408 -2493 434
rect -2644 226 -2493 245
rect -2644 108 -2622 226
rect -2504 108 -2493 226
rect -2644 82 -2493 108
rect -2644 -100 -2493 -81
rect -2644 -218 -2622 -100
rect -2504 -218 -2493 -100
rect -2644 -244 -2493 -218
rect -2644 -426 -2493 -407
rect -2644 -544 -2622 -426
rect -2504 -544 -2493 -426
rect -2644 -570 -2493 -544
rect -2644 -752 -2493 -733
rect -2644 -870 -2622 -752
rect -2504 -870 -2493 -752
rect -2644 -896 -2493 -870
rect -2644 -1079 -2493 -1060
rect -2644 -1197 -2622 -1079
rect -2504 -1197 -2493 -1079
rect -2644 -1223 -2493 -1197
rect -2644 -1406 -2493 -1387
rect -2644 -1524 -2622 -1406
rect -2504 -1524 -2493 -1406
rect -2644 -1550 -2493 -1524
rect -2414 -1511 -2384 3103
rect -2309 2671 -2172 2690
rect -2309 2553 -2294 2671
rect -2176 2553 -2172 2671
rect -2309 2527 -2172 2553
rect -2309 2345 -2172 2364
rect -2309 2227 -2294 2345
rect -2176 2227 -2172 2345
rect -2309 2201 -2172 2227
rect -2309 2019 -2172 2038
rect -2309 1901 -2294 2019
rect -2176 1901 -2172 2019
rect -2309 1875 -2172 1901
rect -2309 1693 -2172 1712
rect -2309 1575 -2294 1693
rect -2176 1575 -2172 1693
rect -2309 1549 -2172 1575
rect -2309 1367 -2172 1386
rect -2309 1249 -2294 1367
rect -2176 1249 -2172 1367
rect -2309 1223 -2172 1249
rect -2092 1194 5604 2862
rect -2092 1187 4143 1194
rect -2092 1069 757 1187
rect 875 1184 4143 1187
rect 875 1069 1059 1184
rect -2092 1066 1059 1069
rect 1177 1161 4143 1184
rect 1177 1066 3847 1161
rect -2309 1041 -2172 1060
rect -2309 923 -2294 1041
rect -2176 923 -2172 1041
rect -2309 897 -2172 923
rect -2092 1043 3847 1066
rect 3965 1076 4143 1161
rect 4261 1076 5604 1194
rect 3965 1043 5604 1076
rect -2309 715 -2172 734
rect -2309 597 -2294 715
rect -2176 597 -2172 715
rect -2309 571 -2172 597
rect -2092 547 5604 1043
rect -2092 540 1040 547
rect -2092 422 767 540
rect 885 429 1040 540
rect 1158 505 5604 547
rect 1158 429 3825 505
rect 885 422 3825 429
rect -2309 389 -2172 408
rect -2309 271 -2294 389
rect -2176 271 -2172 389
rect -2309 245 -2172 271
rect -2092 387 3825 422
rect 3943 488 5604 505
rect 3943 387 4133 488
rect -2092 370 4133 387
rect 4251 370 5604 488
rect -2309 63 -2172 82
rect -2309 -55 -2294 63
rect -2176 -55 -2172 63
rect -2309 -81 -2172 -55
rect -2309 -263 -2172 -244
rect -2309 -381 -2294 -263
rect -2176 -381 -2172 -263
rect -2309 -407 -2172 -381
rect -2309 -589 -2172 -570
rect -2309 -707 -2294 -589
rect -2176 -707 -2172 -589
rect -2309 -733 -2172 -707
rect -2309 -916 -2172 -897
rect -2309 -1034 -2294 -916
rect -2176 -1034 -2172 -916
rect -2309 -1060 -2172 -1034
rect -2092 -1071 5604 370
rect -2092 -1189 -1858 -1071
rect -1740 -1189 5604 -1071
rect -2092 -1250 5604 -1189
rect 851 -1511 894 -1508
rect -2414 -1541 861 -1511
rect 851 -1543 861 -1541
rect 893 -1543 894 -1511
rect 851 -1544 894 -1543
rect 976 -1514 1128 -1512
rect 976 -1515 1091 -1514
rect 976 -1547 977 -1515
rect 1009 -1547 1091 -1515
rect 976 -1548 1091 -1547
rect 1090 -1549 1091 -1548
rect 1127 -1549 1128 -1514
rect 1090 -1550 1128 -1549
rect 1518 -1514 1556 -1513
rect 1518 -1550 1519 -1514
rect 1553 -1515 1668 -1514
rect 1553 -1547 1635 -1515
rect 1667 -1547 1668 -1515
rect 1553 -1550 1668 -1547
rect 1718 -1515 1754 -1250
rect 1718 -1547 1721 -1515
rect 1753 -1547 1754 -1515
rect 1718 -1548 1754 -1547
rect 1863 -1515 1965 -1512
rect 1863 -1547 1864 -1515
rect 1896 -1547 1965 -1515
rect 1863 -1548 1965 -1547
rect 2000 -1548 2010 -1512
rect 2733 -1513 2876 -1512
rect 2404 -1515 2538 -1514
rect 2404 -1549 2405 -1515
rect 2440 -1547 2505 -1515
rect 2537 -1547 2538 -1515
rect 2440 -1549 2538 -1547
rect 2588 -1515 2624 -1513
rect 2588 -1547 2591 -1515
rect 2623 -1547 2624 -1515
rect 2588 -1548 2624 -1547
rect 2733 -1515 2830 -1513
rect 2733 -1547 2734 -1515
rect 2766 -1547 2830 -1515
rect 2864 -1547 2876 -1513
rect 2733 -1548 2876 -1547
rect 3024 -1515 3155 -1514
rect 2404 -1550 2538 -1549
rect 1518 -1551 1556 -1550
rect 2591 -1797 2623 -1548
rect 3024 -1550 3026 -1515
rect 3060 -1547 3122 -1515
rect 3154 -1547 3155 -1515
rect 3060 -1550 3155 -1547
rect 3248 -1515 3298 -1509
rect 3248 -1547 3253 -1515
rect 3285 -1547 3298 -1515
rect 3248 -1797 3298 -1547
rect -2093 -1847 3019 -1797
rect -2093 -1864 725 -1847
rect -2093 -1982 -1843 -1864
rect -1725 -1965 725 -1864
rect 843 -1965 3019 -1847
rect -1725 -1982 3019 -1965
rect -2093 -4825 3019 -1982
rect 3075 -1864 5604 -1797
rect 3075 -1982 3327 -1864
rect 3445 -1982 5604 -1864
rect 3075 -4825 5604 -1982
<< via4 >>
rect -2622 2790 -2504 2834
rect -2622 2758 -2580 2790
rect -2580 2758 -2548 2790
rect -2548 2758 -2504 2790
rect -2622 2716 -2504 2758
rect -2622 2464 -2504 2508
rect -2622 2432 -2580 2464
rect -2580 2432 -2548 2464
rect -2548 2432 -2504 2464
rect -2622 2390 -2504 2432
rect -2622 2138 -2504 2182
rect -2622 2106 -2580 2138
rect -2580 2106 -2548 2138
rect -2548 2106 -2504 2138
rect -2622 2064 -2504 2106
rect -2622 1812 -2504 1856
rect -2622 1780 -2580 1812
rect -2580 1780 -2548 1812
rect -2548 1780 -2504 1812
rect -2622 1738 -2504 1780
rect -2622 1486 -2504 1530
rect -2622 1454 -2580 1486
rect -2580 1454 -2548 1486
rect -2548 1454 -2504 1486
rect -2622 1412 -2504 1454
rect -2622 1160 -2504 1204
rect -2622 1128 -2580 1160
rect -2580 1128 -2548 1160
rect -2548 1128 -2504 1160
rect -2622 1086 -2504 1128
rect -2622 834 -2504 878
rect -2622 802 -2580 834
rect -2580 802 -2548 834
rect -2548 802 -2504 834
rect -2622 760 -2504 802
rect -2622 508 -2504 552
rect -2622 476 -2580 508
rect -2580 476 -2548 508
rect -2548 476 -2504 508
rect -2622 434 -2504 476
rect -2622 182 -2504 226
rect -2622 150 -2580 182
rect -2580 150 -2548 182
rect -2548 150 -2504 182
rect -2622 108 -2504 150
rect -2622 -144 -2504 -100
rect -2622 -176 -2580 -144
rect -2580 -176 -2548 -144
rect -2548 -176 -2504 -144
rect -2622 -218 -2504 -176
rect -2622 -470 -2504 -426
rect -2622 -502 -2580 -470
rect -2580 -502 -2548 -470
rect -2548 -502 -2504 -470
rect -2622 -544 -2504 -502
rect -2622 -796 -2504 -752
rect -2622 -828 -2580 -796
rect -2580 -828 -2548 -796
rect -2548 -828 -2504 -796
rect -2622 -870 -2504 -828
rect -2622 -1123 -2504 -1079
rect -2622 -1155 -2580 -1123
rect -2580 -1155 -2548 -1123
rect -2548 -1155 -2504 -1123
rect -2622 -1197 -2504 -1155
rect -2622 -1450 -2504 -1406
rect -2622 -1482 -2580 -1450
rect -2580 -1482 -2548 -1450
rect -2548 -1482 -2504 -1450
rect -2622 -1524 -2504 -1482
rect -2294 2627 -2176 2671
rect -2294 2595 -2252 2627
rect -2252 2595 -2220 2627
rect -2220 2595 -2176 2627
rect -2294 2553 -2176 2595
rect -2294 2301 -2176 2345
rect -2294 2269 -2252 2301
rect -2252 2269 -2220 2301
rect -2220 2269 -2176 2301
rect -2294 2227 -2176 2269
rect -2294 1975 -2176 2019
rect -2294 1943 -2252 1975
rect -2252 1943 -2220 1975
rect -2220 1943 -2176 1975
rect -2294 1901 -2176 1943
rect -2294 1649 -2176 1693
rect -2294 1617 -2252 1649
rect -2252 1617 -2220 1649
rect -2220 1617 -2176 1649
rect -2294 1575 -2176 1617
rect -2294 1323 -2176 1367
rect -2294 1291 -2252 1323
rect -2252 1291 -2220 1323
rect -2220 1291 -2176 1323
rect -2294 1249 -2176 1291
rect -2294 997 -2176 1041
rect -2294 965 -2252 997
rect -2252 965 -2220 997
rect -2220 965 -2176 997
rect -2294 923 -2176 965
rect -2294 671 -2176 715
rect -2294 639 -2252 671
rect -2252 639 -2220 671
rect -2220 639 -2176 671
rect -2294 597 -2176 639
rect -2294 345 -2176 389
rect -2294 313 -2252 345
rect -2252 313 -2220 345
rect -2220 313 -2176 345
rect -2294 271 -2176 313
rect -2294 19 -2176 63
rect -2294 -13 -2252 19
rect -2252 -13 -2220 19
rect -2220 -13 -2176 19
rect -2294 -55 -2176 -13
rect -2294 -307 -2176 -263
rect -2294 -339 -2252 -307
rect -2252 -339 -2220 -307
rect -2220 -339 -2176 -307
rect -2294 -381 -2176 -339
rect -2294 -633 -2176 -589
rect -2294 -665 -2252 -633
rect -2252 -665 -2220 -633
rect -2220 -665 -2176 -633
rect -2294 -707 -2176 -665
rect -2294 -960 -2176 -916
rect -2294 -992 -2252 -960
rect -2252 -992 -2220 -960
rect -2220 -992 -2176 -960
rect -2294 -1034 -2176 -992
rect 5454 -1575 5572 -1528
rect 5454 -1609 5492 -1575
rect 5492 -1609 5526 -1575
rect 5526 -1609 5572 -1575
rect 5454 -1646 5572 -1609
<< mimcap2 >>
rect -2078 1003 922 2848
rect -2078 885 763 1003
rect 881 885 922 1003
rect -2078 848 922 885
rect 1006 1005 4006 2848
rect 1006 887 1047 1005
rect 1165 987 4006 1005
rect 1165 887 3833 987
rect 1006 869 3833 887
rect 3951 869 4006 987
rect 1006 848 4006 869
rect 4090 992 5590 2848
rect 4090 874 4124 992
rect 4242 874 5590 992
rect 4090 848 5590 874
rect -2078 726 922 764
rect -2078 608 762 726
rect 880 608 922 726
rect -2078 -1089 922 608
rect -2078 -1207 653 -1089
rect 771 -1207 922 -1089
rect -2078 -1236 922 -1207
rect 1006 729 4006 764
rect 1006 611 1044 729
rect 1162 708 4006 729
rect 1162 611 3830 708
rect 1006 590 3830 611
rect 3948 590 4006 708
rect 1006 -1236 4006 590
rect 4090 706 5590 764
rect 4090 588 4122 706
rect 4240 588 5590 706
rect 4090 -1236 5590 588
rect -2079 -1865 421 -1811
rect -2079 -1983 241 -1865
rect 359 -1983 421 -1865
rect -2079 -4811 421 -1983
rect 505 -1865 3005 -1811
rect 505 -1983 554 -1865
rect 672 -1983 3005 -1865
rect 505 -4811 3005 -1983
rect 3089 -1839 5590 -1811
rect 3089 -1957 5450 -1839
rect 5568 -1957 5590 -1839
rect 3089 -4811 5590 -1957
<< mimcap2contact >>
rect 763 885 881 1003
rect 1047 887 1165 1005
rect 3833 869 3951 987
rect 4124 874 4242 992
rect 762 608 880 726
rect 653 -1207 771 -1089
rect 1044 611 1162 729
rect 3830 590 3948 708
rect 4122 588 4240 706
rect 241 -1983 359 -1865
rect 554 -1983 672 -1865
rect 5450 -1957 5568 -1839
<< metal5 >>
rect -2644 2834 -2315 2853
rect -2644 2716 -2622 2834
rect -2504 2716 -2315 2834
rect -2644 2690 -2315 2716
rect -2483 2671 -2155 2690
rect -2483 2553 -2294 2671
rect -2176 2553 -2155 2671
rect -2483 2527 -2155 2553
rect -2644 2508 -2315 2527
rect -2644 2390 -2622 2508
rect -2504 2390 -2315 2508
rect -2644 2364 -2315 2390
rect -2483 2345 -2155 2364
rect -2483 2227 -2294 2345
rect -2176 2227 -2155 2345
rect -2483 2201 -2155 2227
rect -2644 2182 -2315 2201
rect -2644 2064 -2622 2182
rect -2504 2064 -2315 2182
rect -2644 2038 -2315 2064
rect -2483 2019 -2155 2038
rect -2483 1901 -2294 2019
rect -2176 1901 -2155 2019
rect -2483 1875 -2155 1901
rect -2644 1856 -2315 1875
rect -2644 1738 -2622 1856
rect -2504 1738 -2315 1856
rect -2644 1712 -2315 1738
rect -2483 1693 -2155 1712
rect -2483 1575 -2294 1693
rect -2176 1575 -2155 1693
rect -2483 1549 -2155 1575
rect -2644 1530 -2315 1549
rect -2644 1412 -2622 1530
rect -2504 1412 -2315 1530
rect -2644 1386 -2315 1412
rect -2483 1367 -2155 1386
rect -2483 1249 -2294 1367
rect -2176 1249 -2155 1367
rect -2483 1223 -2155 1249
rect -2644 1204 -2315 1223
rect -2644 1086 -2622 1204
rect -2504 1086 -2315 1204
rect -2644 1060 -2315 1086
rect -2483 1041 -2155 1060
rect -2483 923 -2294 1041
rect -2176 923 -2155 1041
rect -2483 897 -2155 923
rect 730 1005 1188 1029
rect 730 1003 1047 1005
rect -2644 878 -2315 897
rect -2644 760 -2622 878
rect -2504 760 -2315 878
rect -2644 734 -2315 760
rect 730 885 763 1003
rect 881 887 1047 1003
rect 1165 887 1188 1005
rect 881 885 1188 887
rect -2483 715 -2155 734
rect -2483 597 -2294 715
rect -2176 597 -2155 715
rect -2483 571 -2155 597
rect 730 729 1188 885
rect 730 726 1044 729
rect 730 608 762 726
rect 880 611 1044 726
rect 1162 611 1188 729
rect 880 608 1188 611
rect 730 592 1188 608
rect 3809 992 4266 1013
rect 3809 987 4124 992
rect 3809 869 3833 987
rect 3951 874 4124 987
rect 4242 874 4266 992
rect 3951 869 4266 874
rect 3809 708 4266 869
rect 3809 590 3830 708
rect 3948 706 4266 708
rect 3948 590 4122 706
rect 3809 588 4122 590
rect 4240 588 4266 706
rect -2644 552 -2315 571
rect 3809 569 4266 588
rect -2644 434 -2622 552
rect -2504 434 -2315 552
rect -2644 408 -2315 434
rect -2483 389 -2155 408
rect -2483 271 -2294 389
rect -2176 271 -2155 389
rect -2483 245 -2155 271
rect -2644 226 -2315 245
rect -2644 108 -2622 226
rect -2504 108 -2315 226
rect -2644 82 -2315 108
rect -2483 63 -2155 82
rect -2483 -55 -2294 63
rect -2176 -55 -2155 63
rect -2483 -81 -2155 -55
rect -2644 -100 -2315 -81
rect -2644 -218 -2622 -100
rect -2504 -218 -2315 -100
rect -2644 -244 -2315 -218
rect -2483 -263 -2155 -244
rect -2483 -381 -2294 -263
rect -2176 -381 -2155 -263
rect -2483 -407 -2155 -381
rect -2644 -426 -2315 -407
rect -2644 -544 -2622 -426
rect -2504 -544 -2315 -426
rect -2644 -570 -2315 -544
rect -2483 -589 -2155 -570
rect -2483 -707 -2294 -589
rect -2176 -707 -2155 -589
rect -2483 -733 -2155 -707
rect -2644 -752 -2315 -733
rect -2644 -870 -2622 -752
rect -2504 -870 -2315 -752
rect -2644 -896 -2315 -870
rect -2483 -897 -2315 -896
rect -2483 -916 -2155 -897
rect -2483 -1034 -2294 -916
rect -2176 -1034 -2155 -916
rect -2483 -1060 -2155 -1034
rect -2644 -1079 -2315 -1060
rect -2644 -1197 -2622 -1079
rect -2504 -1197 -2315 -1079
rect -2644 -1223 -2315 -1197
rect -2483 -1387 -2315 -1223
rect -2644 -1406 -2315 -1387
rect -2644 -1524 -2622 -1406
rect -2504 -1443 -2315 -1406
rect 639 -1089 805 -1073
rect 639 -1207 653 -1089
rect 771 -1207 805 -1089
rect 639 -1443 805 -1207
rect -2504 -1524 839 -1443
rect -2644 -1550 839 -1524
rect -2483 -1609 839 -1550
rect 5428 -1528 5592 -1502
rect 556 -1839 717 -1609
rect 218 -1865 717 -1839
rect 218 -1983 241 -1865
rect 359 -1983 554 -1865
rect 672 -1983 717 -1865
rect 5428 -1646 5454 -1528
rect 5572 -1646 5592 -1528
rect 5428 -1805 5592 -1646
rect 5428 -1839 5591 -1805
rect 5428 -1957 5450 -1839
rect 5568 -1957 5591 -1839
rect 5428 -1978 5591 -1957
rect 218 -2000 717 -1983
<< labels >>
flabel metal4 1885 -36 2909 887 0 FreeSans 800 0 0 0 C1
flabel mimcap 1256 -1622 1447 -1471 0 FreeSans 800 0 0 0 Cs1
rlabel metal4 1033 -1512 1033 -1512 1 cs1
flabel mimcap 2115 -1620 2306 -1469 0 FreeSans 800 0 0 0 Cs2
flabel metal4 -82 -3740 942 -2817 0 FreeSans 800 0 0 0 C2
flabel mimcap2 3912 -3489 4936 -2566 0 FreeSans 800 0 0 0 C3
flabel mimcap 2863 -1593 3054 -1442 0 FreeSans 800 0 0 0 Cs3
rlabel metal4 1754 -1270 1754 -1270 3 c1
rlabel metal4 1922 -1548 1922 -1548 5 cs2
rlabel metal4 2623 -1752 2623 -1752 3 c2
rlabel metal4 3098 -1550 3098 -1550 5 cs3
rlabel metal4 3298 -1734 3298 -1734 3 c3
rlabel metal1 3312 -1741 3312 -1741 3 phi1
rlabel metal1 3313 -1774 3313 -1774 3 phi2
rlabel metal1 3339 -1311 3339 -1311 3 phi1b
rlabel metal1 3337 -1280 3337 -1280 3 phi2b
<< end >>
