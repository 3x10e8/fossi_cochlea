magic
tech sky130A
timestamp 1654156798
use cap_10_10_x2  cap_10_10_x2_0
array 0 3 1098 0 1 1098
timestamp 1654156239
transform 1 0 65 0 1 54
box -57 -52 1041 1046
<< labels >>
flabel space 8 2 4400 2198 0 FreeSans 4000 0 0 0 3.2pF
<< end >>
