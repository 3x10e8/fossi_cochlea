magic
tech sky130B
magscale 1 2
timestamp 1663374946
<< obsli1 >>
rect 1104 2159 406824 21777
<< obsm1 >>
rect 1104 1436 406984 22296
<< metal2 >>
rect 5078 23200 5134 24000
rect 13542 23200 13598 24000
rect 22006 23200 22062 24000
rect 30470 23200 30526 24000
rect 38934 23200 38990 24000
rect 47398 23200 47454 24000
rect 55862 23200 55918 24000
rect 64326 23200 64382 24000
rect 72790 23200 72846 24000
rect 81254 23200 81310 24000
rect 89718 23200 89774 24000
rect 98182 23200 98238 24000
rect 106646 23200 106702 24000
rect 115110 23200 115166 24000
rect 123574 23200 123630 24000
rect 132038 23200 132094 24000
rect 140502 23200 140558 24000
rect 148966 23200 149022 24000
rect 157430 23200 157486 24000
rect 165894 23200 165950 24000
rect 174358 23200 174414 24000
rect 182822 23200 182878 24000
rect 191286 23200 191342 24000
rect 199750 23200 199806 24000
rect 208214 23200 208270 24000
rect 216678 23200 216734 24000
rect 225142 23200 225198 24000
rect 233606 23200 233662 24000
rect 242070 23200 242126 24000
rect 250534 23200 250590 24000
rect 258998 23200 259054 24000
rect 267462 23200 267518 24000
rect 275926 23200 275982 24000
rect 284390 23200 284446 24000
rect 292854 23200 292910 24000
rect 301318 23200 301374 24000
rect 309782 23200 309838 24000
rect 318246 23200 318302 24000
rect 326710 23200 326766 24000
rect 335174 23200 335230 24000
rect 343638 23200 343694 24000
rect 352102 23200 352158 24000
rect 360566 23200 360622 24000
rect 369030 23200 369086 24000
rect 377494 23200 377550 24000
rect 385958 23200 386014 24000
rect 394422 23200 394478 24000
rect 402886 23200 402942 24000
rect 5078 0 5134 800
rect 13542 0 13598 800
rect 22006 0 22062 800
rect 30470 0 30526 800
rect 38934 0 38990 800
rect 47398 0 47454 800
rect 55862 0 55918 800
rect 64326 0 64382 800
rect 72790 0 72846 800
rect 81254 0 81310 800
rect 89718 0 89774 800
rect 98182 0 98238 800
rect 106646 0 106702 800
rect 115110 0 115166 800
rect 123574 0 123630 800
rect 132038 0 132094 800
rect 140502 0 140558 800
rect 148966 0 149022 800
rect 157430 0 157486 800
rect 165894 0 165950 800
rect 174358 0 174414 800
rect 182822 0 182878 800
rect 191286 0 191342 800
rect 199750 0 199806 800
rect 208214 0 208270 800
rect 216678 0 216734 800
rect 225142 0 225198 800
rect 233606 0 233662 800
rect 242070 0 242126 800
rect 250534 0 250590 800
rect 258998 0 259054 800
rect 267462 0 267518 800
rect 275926 0 275982 800
rect 284390 0 284446 800
rect 292854 0 292910 800
rect 301318 0 301374 800
rect 309782 0 309838 800
rect 318246 0 318302 800
rect 326710 0 326766 800
rect 335174 0 335230 800
rect 343638 0 343694 800
rect 352102 0 352158 800
rect 360566 0 360622 800
rect 369030 0 369086 800
rect 377494 0 377550 800
rect 385958 0 386014 800
rect 394422 0 394478 800
rect 402886 0 402942 800
<< obsm2 >>
rect 1582 23144 5022 23338
rect 5190 23144 13486 23338
rect 13654 23144 21950 23338
rect 22118 23144 30414 23338
rect 30582 23144 38878 23338
rect 39046 23144 47342 23338
rect 47510 23144 55806 23338
rect 55974 23144 64270 23338
rect 64438 23144 72734 23338
rect 72902 23144 81198 23338
rect 81366 23144 89662 23338
rect 89830 23144 98126 23338
rect 98294 23144 106590 23338
rect 106758 23144 115054 23338
rect 115222 23144 123518 23338
rect 123686 23144 131982 23338
rect 132150 23144 140446 23338
rect 140614 23144 148910 23338
rect 149078 23144 157374 23338
rect 157542 23144 165838 23338
rect 166006 23144 174302 23338
rect 174470 23144 182766 23338
rect 182934 23144 191230 23338
rect 191398 23144 199694 23338
rect 199862 23144 208158 23338
rect 208326 23144 216622 23338
rect 216790 23144 225086 23338
rect 225254 23144 233550 23338
rect 233718 23144 242014 23338
rect 242182 23144 250478 23338
rect 250646 23144 258942 23338
rect 259110 23144 267406 23338
rect 267574 23144 275870 23338
rect 276038 23144 284334 23338
rect 284502 23144 292798 23338
rect 292966 23144 301262 23338
rect 301430 23144 309726 23338
rect 309894 23144 318190 23338
rect 318358 23144 326654 23338
rect 326822 23144 335118 23338
rect 335286 23144 343582 23338
rect 343750 23144 352046 23338
rect 352214 23144 360510 23338
rect 360678 23144 368974 23338
rect 369142 23144 377438 23338
rect 377606 23144 385902 23338
rect 386070 23144 394366 23338
rect 394534 23144 402830 23338
rect 402998 23144 406978 23338
rect 1582 856 406978 23144
rect 1582 734 5022 856
rect 5190 734 13486 856
rect 13654 734 21950 856
rect 22118 734 30414 856
rect 30582 734 38878 856
rect 39046 734 47342 856
rect 47510 734 55806 856
rect 55974 734 64270 856
rect 64438 734 72734 856
rect 72902 734 81198 856
rect 81366 734 89662 856
rect 89830 734 98126 856
rect 98294 734 106590 856
rect 106758 734 115054 856
rect 115222 734 123518 856
rect 123686 734 131982 856
rect 132150 734 140446 856
rect 140614 734 148910 856
rect 149078 734 157374 856
rect 157542 734 165838 856
rect 166006 734 174302 856
rect 174470 734 182766 856
rect 182934 734 191230 856
rect 191398 734 199694 856
rect 199862 734 208158 856
rect 208326 734 216622 856
rect 216790 734 225086 856
rect 225254 734 233550 856
rect 233718 734 242014 856
rect 242182 734 250478 856
rect 250646 734 258942 856
rect 259110 734 267406 856
rect 267574 734 275870 856
rect 276038 734 284334 856
rect 284502 734 292798 856
rect 292966 734 301262 856
rect 301430 734 309726 856
rect 309894 734 318190 856
rect 318358 734 326654 856
rect 326822 734 335118 856
rect 335286 734 343582 856
rect 343750 734 352046 856
rect 352214 734 360510 856
rect 360678 734 368974 856
rect 369142 734 377438 856
rect 377606 734 385902 856
rect 386070 734 394366 856
rect 394534 734 402830 856
rect 402998 734 406978 856
<< metal3 >>
rect 0 22040 800 22160
rect 0 18640 800 18760
rect 0 15240 800 15360
rect 0 11840 800 11960
rect 0 8440 800 8560
rect 0 5040 800 5160
rect 0 1640 800 1760
<< obsm3 >>
rect 800 22240 406982 22269
rect 880 21960 406982 22240
rect 800 18840 406982 21960
rect 880 18560 406982 18840
rect 800 15440 406982 18560
rect 880 15160 406982 15440
rect 800 12040 406982 15160
rect 880 11760 406982 12040
rect 800 8640 406982 11760
rect 880 8360 406982 8640
rect 800 5240 406982 8360
rect 880 4960 406982 5240
rect 800 1840 406982 4960
rect 880 1667 406982 1840
<< metal4 >>
rect 51659 2128 51979 21808
rect 102374 2128 102694 21808
rect 153089 2128 153409 21808
rect 203804 2128 204124 21808
rect 254519 2128 254839 21808
rect 305234 2128 305554 21808
rect 355949 2128 356269 21808
rect 406664 2128 406984 21808
<< obsm4 >>
rect 9075 21888 403085 22269
rect 9075 2483 51579 21888
rect 52059 2483 102294 21888
rect 102774 2483 153009 21888
rect 153489 2483 203724 21888
rect 204204 2483 254439 21888
rect 254919 2483 305154 21888
rect 305634 2483 355869 21888
rect 356349 2483 403085 21888
<< labels >>
rlabel metal2 s 13542 23200 13598 24000 6 cclk_I[0]
port 1 nsew signal output
rlabel metal2 s 64326 23200 64382 24000 6 cclk_I[1]
port 2 nsew signal output
rlabel metal2 s 115110 23200 115166 24000 6 cclk_I[2]
port 3 nsew signal output
rlabel metal2 s 165894 23200 165950 24000 6 cclk_I[3]
port 4 nsew signal output
rlabel metal2 s 216678 23200 216734 24000 6 cclk_I[4]
port 5 nsew signal output
rlabel metal2 s 267462 23200 267518 24000 6 cclk_I[5]
port 6 nsew signal output
rlabel metal2 s 318246 23200 318302 24000 6 cclk_I[6]
port 7 nsew signal output
rlabel metal2 s 369030 23200 369086 24000 6 cclk_I[7]
port 8 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 cclk_Q[0]
port 9 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 cclk_Q[1]
port 10 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 cclk_Q[2]
port 11 nsew signal output
rlabel metal2 s 165894 0 165950 800 6 cclk_Q[3]
port 12 nsew signal output
rlabel metal2 s 216678 0 216734 800 6 cclk_Q[4]
port 13 nsew signal output
rlabel metal2 s 267462 0 267518 800 6 cclk_Q[5]
port 14 nsew signal output
rlabel metal2 s 318246 0 318302 800 6 cclk_Q[6]
port 15 nsew signal output
rlabel metal2 s 369030 0 369086 800 6 cclk_Q[7]
port 16 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 clk_master
port 17 nsew signal input
rlabel metal2 s 22006 23200 22062 24000 6 clkdiv2_I[0]
port 18 nsew signal output
rlabel metal2 s 72790 23200 72846 24000 6 clkdiv2_I[1]
port 19 nsew signal output
rlabel metal2 s 123574 23200 123630 24000 6 clkdiv2_I[2]
port 20 nsew signal output
rlabel metal2 s 174358 23200 174414 24000 6 clkdiv2_I[3]
port 21 nsew signal output
rlabel metal2 s 225142 23200 225198 24000 6 clkdiv2_I[4]
port 22 nsew signal output
rlabel metal2 s 275926 23200 275982 24000 6 clkdiv2_I[5]
port 23 nsew signal output
rlabel metal2 s 326710 23200 326766 24000 6 clkdiv2_I[6]
port 24 nsew signal output
rlabel metal2 s 377494 23200 377550 24000 6 clkdiv2_I[7]
port 25 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 clkdiv2_Q[0]
port 26 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 clkdiv2_Q[1]
port 27 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 clkdiv2_Q[2]
port 28 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 clkdiv2_Q[3]
port 29 nsew signal output
rlabel metal2 s 225142 0 225198 800 6 clkdiv2_Q[4]
port 30 nsew signal output
rlabel metal2 s 275926 0 275982 800 6 clkdiv2_Q[5]
port 31 nsew signal output
rlabel metal2 s 326710 0 326766 800 6 clkdiv2_Q[6]
port 32 nsew signal output
rlabel metal2 s 377494 0 377550 800 6 clkdiv2_Q[7]
port 33 nsew signal output
rlabel metal2 s 30470 23200 30526 24000 6 comp_high_I[0]
port 34 nsew signal input
rlabel metal2 s 81254 23200 81310 24000 6 comp_high_I[1]
port 35 nsew signal input
rlabel metal2 s 132038 23200 132094 24000 6 comp_high_I[2]
port 36 nsew signal input
rlabel metal2 s 182822 23200 182878 24000 6 comp_high_I[3]
port 37 nsew signal input
rlabel metal2 s 233606 23200 233662 24000 6 comp_high_I[4]
port 38 nsew signal input
rlabel metal2 s 284390 23200 284446 24000 6 comp_high_I[5]
port 39 nsew signal input
rlabel metal2 s 335174 23200 335230 24000 6 comp_high_I[6]
port 40 nsew signal input
rlabel metal2 s 385958 23200 386014 24000 6 comp_high_I[7]
port 41 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 comp_high_Q[0]
port 42 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 comp_high_Q[1]
port 43 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 comp_high_Q[2]
port 44 nsew signal input
rlabel metal2 s 182822 0 182878 800 6 comp_high_Q[3]
port 45 nsew signal input
rlabel metal2 s 233606 0 233662 800 6 comp_high_Q[4]
port 46 nsew signal input
rlabel metal2 s 284390 0 284446 800 6 comp_high_Q[5]
port 47 nsew signal input
rlabel metal2 s 335174 0 335230 800 6 comp_high_Q[6]
port 48 nsew signal input
rlabel metal2 s 385958 0 386014 800 6 comp_high_Q[7]
port 49 nsew signal input
rlabel metal2 s 47398 23200 47454 24000 6 cos_out[0]
port 50 nsew signal output
rlabel metal2 s 98182 23200 98238 24000 6 cos_out[1]
port 51 nsew signal output
rlabel metal2 s 148966 23200 149022 24000 6 cos_out[2]
port 52 nsew signal output
rlabel metal2 s 199750 23200 199806 24000 6 cos_out[3]
port 53 nsew signal output
rlabel metal2 s 250534 23200 250590 24000 6 cos_out[4]
port 54 nsew signal output
rlabel metal2 s 301318 23200 301374 24000 6 cos_out[5]
port 55 nsew signal output
rlabel metal2 s 352102 23200 352158 24000 6 cos_out[6]
port 56 nsew signal output
rlabel metal2 s 402886 23200 402942 24000 6 cos_out[7]
port 57 nsew signal output
rlabel metal2 s 5078 23200 5134 24000 6 fb1_I[0]
port 58 nsew signal output
rlabel metal2 s 55862 23200 55918 24000 6 fb1_I[1]
port 59 nsew signal output
rlabel metal2 s 106646 23200 106702 24000 6 fb1_I[2]
port 60 nsew signal output
rlabel metal2 s 157430 23200 157486 24000 6 fb1_I[3]
port 61 nsew signal output
rlabel metal2 s 208214 23200 208270 24000 6 fb1_I[4]
port 62 nsew signal output
rlabel metal2 s 258998 23200 259054 24000 6 fb1_I[5]
port 63 nsew signal output
rlabel metal2 s 309782 23200 309838 24000 6 fb1_I[6]
port 64 nsew signal output
rlabel metal2 s 360566 23200 360622 24000 6 fb1_I[7]
port 65 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 fb1_Q[0]
port 66 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 fb1_Q[1]
port 67 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 fb1_Q[2]
port 68 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 fb1_Q[3]
port 69 nsew signal output
rlabel metal2 s 208214 0 208270 800 6 fb1_Q[4]
port 70 nsew signal output
rlabel metal2 s 258998 0 259054 800 6 fb1_Q[5]
port 71 nsew signal output
rlabel metal2 s 309782 0 309838 800 6 fb1_Q[6]
port 72 nsew signal output
rlabel metal2 s 360566 0 360622 800 6 fb1_Q[7]
port 73 nsew signal output
rlabel metal2 s 38934 23200 38990 24000 6 phi1b_dig_I[0]
port 74 nsew signal input
rlabel metal2 s 89718 23200 89774 24000 6 phi1b_dig_I[1]
port 75 nsew signal input
rlabel metal2 s 140502 23200 140558 24000 6 phi1b_dig_I[2]
port 76 nsew signal input
rlabel metal2 s 191286 23200 191342 24000 6 phi1b_dig_I[3]
port 77 nsew signal input
rlabel metal2 s 242070 23200 242126 24000 6 phi1b_dig_I[4]
port 78 nsew signal input
rlabel metal2 s 292854 23200 292910 24000 6 phi1b_dig_I[5]
port 79 nsew signal input
rlabel metal2 s 343638 23200 343694 24000 6 phi1b_dig_I[6]
port 80 nsew signal input
rlabel metal2 s 394422 23200 394478 24000 6 phi1b_dig_I[7]
port 81 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 phi1b_dig_Q[0]
port 82 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 phi1b_dig_Q[1]
port 83 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 phi1b_dig_Q[2]
port 84 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 phi1b_dig_Q[3]
port 85 nsew signal input
rlabel metal2 s 242070 0 242126 800 6 phi1b_dig_Q[4]
port 86 nsew signal input
rlabel metal2 s 292854 0 292910 800 6 phi1b_dig_Q[5]
port 87 nsew signal input
rlabel metal2 s 343638 0 343694 800 6 phi1b_dig_Q[6]
port 88 nsew signal input
rlabel metal2 s 394422 0 394478 800 6 phi1b_dig_Q[7]
port 89 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 read_out_I[0]
port 90 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 read_out_I[1]
port 91 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 read_out_Q[0]
port 92 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 read_out_Q[1]
port 93 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 rstb
port 94 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 sin_out[0]
port 95 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 sin_out[1]
port 96 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 sin_out[2]
port 97 nsew signal output
rlabel metal2 s 199750 0 199806 800 6 sin_out[3]
port 98 nsew signal output
rlabel metal2 s 250534 0 250590 800 6 sin_out[4]
port 99 nsew signal output
rlabel metal2 s 301318 0 301374 800 6 sin_out[5]
port 100 nsew signal output
rlabel metal2 s 352102 0 352158 800 6 sin_out[6]
port 101 nsew signal output
rlabel metal2 s 402886 0 402942 800 6 sin_out[7]
port 102 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 ud_en
port 103 nsew signal input
rlabel metal4 s 51659 2128 51979 21808 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 153089 2128 153409 21808 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 254519 2128 254839 21808 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 355949 2128 356269 21808 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 102374 2128 102694 21808 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 203804 2128 204124 21808 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 305234 2128 305554 21808 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 406664 2128 406984 21808 6 vssd1
port 105 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 408000 24000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14610318
string GDS_FILE /local_disk/fossi_cochlea/openlane/digital_unison/runs/22_09_16_17_31/results/signoff/digital_unison.magic.gds
string GDS_START 632598
<< end >>

