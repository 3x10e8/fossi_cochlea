magic
tech sky130B
magscale 1 2
timestamp 1654741520
use cap_10_10__side_x2  cap_10_10__side_x2_0
array 0 0 -3056 0 5 2720
timestamp 1654741520
transform 0 1 748 -1 0 2727
box -712 -366 2344 2354
use cap_10_10__side_x2  cap_10_10__side_x2_1
array 0 0 -3056 0 5 2720
timestamp 1654741520
transform 0 -1 16336 1 0 -1961
box -712 -366 2344 2354
use cap_10_10_edge_x2  cap_10_10_edge_x2_0
timestamp 1654741520
transform 1 0 -1962 0 1 -1971
box -712 -702 2344 2354
use cap_10_10_edge_x2  cap_10_10_edge_x2_1
timestamp 1654741520
transform 0 1 -1972 -1 0 2727
box -712 -702 2344 2354
use cap_10_10_edge_x2  cap_10_10_edge_x2_2
timestamp 1654741520
transform 0 -1 19056 1 0 -1961
box -712 -702 2344 2354
use cap_10_10_edge_x2  cap_10_10_edge_x2_3
timestamp 1654741520
transform -1 0 19046 0 -1 2737
box -712 -702 2344 2354
<< end >>
