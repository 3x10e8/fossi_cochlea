magic
tech sky130A
magscale 1 2
timestamp 1654311152
<< metal2 >>
rect -10241 27926 -10232 27982
rect -10176 27926 -10167 27982
rect -8477 27925 -8468 27981
rect -8412 27925 -8403 27981
rect 1569 27738 1626 27747
rect 1569 27673 1626 27682
rect 2994 27738 3050 27747
rect 2994 27673 3050 27682
rect 8509 27596 8565 27605
rect 8509 27531 8565 27540
rect 9535 27596 9591 27605
rect 9535 27531 9591 27540
<< via2 >>
rect -10232 27926 -10176 27982
rect -8468 27925 -8412 27981
rect 1569 27682 1626 27738
rect 2994 27682 3050 27738
rect 8509 27540 8565 27596
rect 9535 27540 9591 27596
<< metal3 >>
rect -10241 27982 -9936 27987
rect -10241 27926 -10232 27982
rect -10176 27926 -9936 27982
rect -10241 27921 -9936 27926
rect -8710 27981 -8402 27986
rect -8710 27925 -8468 27981
rect -8412 27925 -8402 27981
rect -8710 27920 -8402 27925
rect 1564 27738 1789 27743
rect 1564 27682 1569 27738
rect 1626 27682 1789 27738
rect 1564 27677 1789 27682
rect 2830 27738 3055 27743
rect 2830 27682 2994 27738
rect 3050 27682 3055 27738
rect 2830 27677 3055 27682
rect 8504 27596 8728 27601
rect 8504 27540 8509 27596
rect 8565 27540 8728 27596
rect 8504 27535 8728 27540
rect 9371 27596 9596 27601
rect 9371 27540 9535 27596
rect 9591 27540 9596 27596
rect 9371 27535 9596 27540
rect -9711 27215 -9529 27517
rect 2242 27044 2344 27504
rect 8978 27201 9110 27515
rect 8323 27112 9110 27201
rect 1370 26963 2344 27044
rect 1351 26279 2784 26410
rect 1351 26215 2113 26279
rect 2177 26215 2784 26279
rect 1351 26090 2784 26215
rect 1362 22673 2795 22810
rect 1362 22609 2110 22673
rect 2174 22609 2795 22673
rect 1362 22490 2795 22609
rect 1369 19219 2802 19332
rect 1369 19155 2133 19219
rect 2197 19155 2802 19219
rect 1369 19012 2802 19155
rect 1360 15745 2793 15879
rect 1360 15681 2095 15745
rect 2159 15681 2793 15745
rect 1360 15559 2793 15681
rect 1367 12259 2800 12381
rect 1367 12195 2102 12259
rect 2166 12195 2800 12259
rect 1367 12061 2800 12195
rect 1373 8771 2806 8906
rect 1373 8707 2073 8771
rect 2137 8707 2806 8771
rect 1373 8586 2806 8707
rect 1365 5322 2798 5457
rect 1365 5258 2075 5322
rect 2139 5258 2798 5322
rect 1365 5137 2798 5258
rect 1358 1817 2791 1935
rect 1358 1753 2055 1817
rect 2119 1753 2791 1817
rect 1358 1615 2791 1753
<< via3 >>
rect 2113 26215 2177 26279
rect 2110 22609 2174 22673
rect 2133 19155 2197 19219
rect 2095 15681 2159 15745
rect 2102 12195 2166 12259
rect 2073 8707 2137 8771
rect 2075 5258 2139 5322
rect 2055 1753 2119 1817
<< metal4 >>
rect -10135 28126 -9830 28198
rect -8751 28126 -8490 28198
rect -8137 28126 -8023 28198
rect -8083 27118 -8023 28126
rect 1126 27890 1298 27962
rect 1688 27890 1786 27962
rect 2832 27890 2930 27962
rect 3316 27896 3394 27962
rect 1126 27212 1286 27890
rect 3262 27811 3394 27896
rect 3316 27193 3394 27811
rect 8089 27749 8249 27820
rect 8089 27669 8313 27749
rect 8636 27748 8734 27820
rect 9370 27748 9468 27820
rect 9832 27751 9992 27820
rect 9802 27669 9992 27751
rect 8089 27228 8249 27669
rect 9832 27226 9992 27669
rect 2024 26367 2277 26368
rect 2024 26131 2032 26367
rect 2268 26131 2277 26367
rect 2021 22761 2274 22762
rect 2021 22525 2029 22761
rect 2265 22525 2274 22761
rect 2044 19307 2297 19308
rect 2044 19071 2052 19307
rect 2288 19071 2297 19307
rect 2006 15833 2259 15834
rect 2006 15597 2014 15833
rect 2250 15597 2259 15833
rect 2013 12347 2266 12348
rect 2013 12111 2021 12347
rect 2257 12111 2266 12347
rect 1984 8859 2237 8860
rect 1984 8623 1992 8859
rect 2228 8623 2237 8859
rect 1986 5410 2239 5411
rect 1986 5174 1994 5410
rect 2230 5174 2239 5410
rect 1966 1905 2219 1906
rect 1966 1669 1974 1905
rect 2210 1669 2219 1905
<< via4 >>
rect 2032 26279 2268 26367
rect 2032 26215 2113 26279
rect 2113 26215 2177 26279
rect 2177 26215 2268 26279
rect 2032 26131 2268 26215
rect 2029 22673 2265 22761
rect 2029 22609 2110 22673
rect 2110 22609 2174 22673
rect 2174 22609 2265 22673
rect 2029 22525 2265 22609
rect 2052 19219 2288 19307
rect 2052 19155 2133 19219
rect 2133 19155 2197 19219
rect 2197 19155 2288 19219
rect 2052 19071 2288 19155
rect 2014 15745 2250 15833
rect 2014 15681 2095 15745
rect 2095 15681 2159 15745
rect 2159 15681 2250 15745
rect 2014 15597 2250 15681
rect 2021 12259 2257 12347
rect 2021 12195 2102 12259
rect 2102 12195 2166 12259
rect 2166 12195 2257 12259
rect 2021 12111 2257 12195
rect 1992 8771 2228 8859
rect 1992 8707 2073 8771
rect 2073 8707 2137 8771
rect 2137 8707 2228 8771
rect 1992 8623 2228 8707
rect 1994 5322 2230 5410
rect 1994 5258 2075 5322
rect 2075 5258 2139 5322
rect 2139 5258 2230 5322
rect 1994 5174 2230 5258
rect 1974 1817 2210 1905
rect 1974 1753 2055 1817
rect 2055 1753 2119 1817
rect 2119 1753 2210 1817
rect 1974 1669 2210 1753
<< metal5 >>
rect 1351 26367 2784 26410
rect 1351 26131 2032 26367
rect 2268 26131 2784 26367
rect 1351 26090 2784 26131
rect 1362 22761 2795 22810
rect 1362 22525 2029 22761
rect 2265 22525 2795 22761
rect 1362 22490 2795 22525
rect 1369 19307 2802 19332
rect 1369 19071 2052 19307
rect 2288 19071 2802 19307
rect 1369 19012 2802 19071
rect 1360 15833 2793 15879
rect 1360 15597 2014 15833
rect 2250 15597 2793 15833
rect 1360 15559 2793 15597
rect 1367 12347 2800 12381
rect 1367 12111 2021 12347
rect 2257 12111 2800 12347
rect 1367 12061 2800 12111
rect 1373 8859 2806 8906
rect 1373 8623 1992 8859
rect 2228 8623 2806 8859
rect 1373 8586 2806 8623
rect 1365 5410 2798 5457
rect 1365 5174 1994 5410
rect 2230 5174 2798 5410
rect 1365 5137 2798 5174
rect 1358 1905 2791 1935
rect 1358 1669 1974 1905
rect 2210 1669 2791 1905
rect 1358 1615 2791 1669
use cap_3pF_8x1  cap_3pF_8x1_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 0 -1 11832 1 0 3532
box -2794 0 23698 2104
use cap_6pF_8x2  cap_6pF_8x2_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 0 -1 8353 1 0 3532
box -2794 0 23698 5588
use cap_10fF  cap_10fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 0 -1 9349 1 0 27529
box -28 -28 708 628
use cap_12pF  cap_12pF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 0 -1 -1404 1 0 3558
box -2820 -2794 23672 9762
use cap_20fF  cap_20fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 0 -1 2809 1 0 27514
box -28 -28 828 1028
use cap_40fF  cap_40fF_0 ~/Documents/fossi_cochlea/mag/final_designs/caps
timestamp 1654307754
transform 0 -1 -8732 1 0 27498
box -28 -28 1368 1228
use cmos_switch_fin  cmos_switch_0 ./filter
timestamp 1654308691
transform 1 0 -10337 0 1 28009
box -175 -95 235 381
use cmos_switch_fin  cmos_switch_1
timestamp 1654308691
transform -1 0 -8307 0 1 28009
box -175 -95 235 381
use cmos_switch_fin  cmos_switch_2
timestamp 1654308691
transform 1 0 1465 0 1 27773
box -175 -95 235 381
use cmos_switch_fin  cmos_switch_3
timestamp 1654308691
transform -1 0 3154 0 1 27773
box -175 -95 235 381
use cmos_switch_fin  cmos_switch_4
timestamp 1654308691
transform 1 0 8405 0 1 27631
box -175 -95 235 381
use cmos_switch_fin  cmos_switch_5
timestamp 1654308691
transform -1 0 9695 0 1 27631
box -175 -95 235 381
<< end >>
