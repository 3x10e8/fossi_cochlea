magic
tech sky130A
magscale 1 2
timestamp 1647910990
<< error_s >>
rect 8765 14234 8771 14240
rect 11557 14234 11563 14240
rect 3754 14225 3774 14231
rect 6146 14225 6166 14231
rect 8797 14210 8801 14230
rect 11527 14210 11531 14230
rect 4299 14199 4308 14209
rect 6691 14199 6700 14209
rect 7511 14207 7524 14209
rect 7558 14207 7577 14209
rect 7558 14199 7559 14207
rect 3732 14177 3733 14189
rect 6124 14177 6125 14189
rect 4265 14165 4274 14175
rect 6657 14165 6666 14175
rect 7477 14173 7490 14175
rect 7592 14173 7611 14175
rect 7592 14165 7593 14173
rect 3703 14147 3715 14159
rect 6095 14147 6107 14159
rect 3971 14126 3983 14135
rect 6363 14126 6375 14135
rect 8839 14122 8843 14142
rect 11485 14122 11489 14142
rect 8795 14100 8801 14106
rect 11527 14100 11533 14106
rect 4009 14088 4021 14097
rect 6401 14088 6413 14097
rect 3147 14073 3164 14079
rect 5539 14073 5556 14079
rect 2509 13744 2515 13750
rect 3403 13744 3420 13745
rect 2541 13720 2545 13740
rect 3437 13710 3454 13711
rect 2583 13632 2587 13652
rect 8421 13645 8437 13647
rect 10053 13645 10066 13647
rect 10168 13645 10187 13647
rect 2539 13610 2545 13616
rect 8387 13611 8403 13613
rect 10087 13611 10100 13613
rect 10134 13611 10153 13613
rect 3371 13119 3384 13121
rect 3418 13119 3437 13121
rect 6407 13119 6420 13121
rect 6454 13119 6473 13121
rect 7783 13119 7802 13121
rect 7836 13119 7849 13121
rect 9347 13119 9366 13121
rect 9400 13119 9413 13121
rect 11331 13119 11347 13121
rect 3418 13111 3419 13119
rect 3337 13085 3350 13087
rect 3452 13085 3471 13087
rect 6373 13085 6386 13087
rect 6488 13085 6507 13087
rect 7749 13085 7768 13087
rect 7870 13085 7883 13087
rect 9313 13085 9332 13087
rect 9434 13085 9447 13087
rect 11365 13085 11381 13087
rect 3452 13077 3453 13085
rect 11741 12656 11747 12662
rect 3050 12635 3051 12641
rect 11711 12632 11715 12652
rect 3084 12601 3085 12607
rect 7675 12559 7676 12567
rect 2969 12557 2982 12559
rect 3084 12557 3103 12559
rect 4465 12557 4481 12559
rect 5913 12557 5926 12559
rect 6028 12557 6047 12559
rect 7657 12557 7676 12559
rect 7778 12557 7791 12559
rect 8303 12557 8319 12559
rect 10329 12557 10342 12559
rect 10444 12557 10463 12559
rect 10971 12557 10987 12559
rect 11669 12544 11673 12564
rect 7709 12525 7710 12533
rect 3003 12523 3016 12525
rect 3050 12523 3069 12525
rect 4431 12523 4447 12525
rect 5947 12523 5960 12525
rect 5994 12523 6013 12525
rect 7691 12523 7710 12525
rect 7744 12523 7757 12525
rect 8337 12523 8353 12525
rect 10363 12523 10376 12525
rect 10410 12523 10429 12525
rect 11005 12523 11021 12525
rect 11711 12522 11717 12528
rect 3723 12230 3732 12236
rect 3695 12202 3704 12208
rect 2509 12058 2515 12064
rect 2541 12034 2545 12054
rect 5487 12031 5500 12033
rect 5534 12031 5553 12033
rect 5453 11997 5466 11999
rect 5568 11997 5587 11999
rect 2583 11946 2587 11966
rect 2539 11924 2545 11930
rect 11146 11603 11163 11609
rect 10327 11547 10339 11556
rect 10675 11527 10687 11539
rect 10365 11509 10377 11518
rect 10645 11485 10646 11497
rect 3085 11469 3101 11471
rect 5083 11469 5099 11471
rect 6369 11469 6388 11471
rect 6490 11469 6503 11471
rect 10074 11469 10083 11479
rect 10616 11455 10636 11461
rect 3051 11435 3067 11437
rect 5117 11435 5133 11437
rect 6403 11435 6422 11437
rect 6456 11435 6469 11437
rect 10040 11435 10049 11445
rect 10892 11142 10900 11148
rect 10920 11114 10928 11120
rect 3122 10961 3142 10967
rect 2588 10935 2597 10945
rect 7191 10943 7207 10945
rect 7835 10943 7851 10945
rect 8891 10943 8904 10945
rect 8938 10943 8957 10945
rect 10451 10943 10470 10945
rect 10504 10943 10517 10945
rect 3163 10913 3164 10925
rect 2622 10901 2631 10911
rect 7225 10909 7241 10911
rect 7869 10909 7885 10911
rect 8857 10909 8870 10911
rect 8972 10909 8991 10911
rect 10417 10909 10436 10911
rect 10538 10909 10551 10911
rect 3181 10883 3193 10895
rect 2913 10862 2925 10871
rect 2875 10824 2887 10833
rect 3732 10809 3749 10815
rect 3829 10515 3846 10521
rect 9398 10515 9415 10521
rect 2509 10480 2515 10486
rect 6129 10480 6135 10486
rect 10637 10480 10643 10486
rect 11617 10480 11623 10486
rect 2541 10456 2545 10476
rect 4653 10459 4665 10468
rect 6099 10456 6103 10476
rect 8579 10459 8591 10468
rect 10607 10456 10611 10476
rect 11649 10456 11653 10476
rect 4305 10439 4317 10451
rect 8927 10439 8939 10451
rect 4615 10421 4627 10430
rect 8617 10421 8629 10430
rect 4346 10397 4347 10409
rect 8897 10397 8898 10409
rect 2583 10368 2587 10388
rect 4909 10381 4918 10391
rect 4356 10367 4376 10373
rect 6057 10368 6061 10388
rect 8326 10381 8335 10391
rect 8868 10367 8888 10373
rect 10565 10368 10569 10388
rect 11691 10368 11695 10388
rect 2539 10346 2545 10352
rect 4943 10347 4952 10357
rect 6099 10346 6105 10352
rect 8292 10347 8301 10357
rect 10607 10346 10613 10352
rect 11647 10346 11653 10352
rect 6238 9873 6258 9879
rect 11206 9873 11226 9879
rect 6783 9847 6792 9857
rect 8797 9855 8813 9857
rect 11751 9847 11760 9857
rect 6216 9825 6217 9837
rect 11184 9825 11185 9837
rect 6749 9813 6758 9823
rect 8763 9821 8779 9823
rect 11717 9813 11726 9823
rect 6187 9795 6199 9807
rect 11155 9795 11167 9807
rect 6455 9774 6467 9783
rect 11423 9774 11435 9783
rect 3534 9757 3551 9758
rect 6493 9736 6505 9745
rect 11461 9736 11473 9745
rect 3568 9723 3585 9724
rect 5631 9721 5648 9727
rect 10599 9721 10616 9727
<< nwell >>
rect 14580 11851 14755 12005
<< locali >>
rect 14927 11592 14959 11593
rect 14927 11462 14961 11592
<< viali >>
rect 14926 11764 14961 11800
rect 15036 11721 15070 11755
rect 14926 11677 14960 11711
rect 14547 11543 14583 11579
rect 15037 11384 15071 11418
rect 14927 11340 14961 11374
rect 14927 11252 14961 11286
rect 14549 11206 14583 11240
<< metal1 >>
rect 16975 13103 17027 13109
rect 16568 13061 16975 13095
rect 16975 13045 17027 13051
rect 17185 12728 17237 12734
rect 16544 12681 17185 12715
rect 17185 12665 17237 12671
rect 17115 12474 17167 12480
rect 15002 12421 15008 12473
rect 15060 12421 15066 12473
rect 16544 12429 17115 12463
rect 17115 12409 17167 12415
rect 14533 12103 14595 12110
rect 16906 12093 16958 12099
rect 16575 12049 16906 12083
rect 14533 12028 14595 12035
rect 16906 12033 16958 12039
rect 14898 11752 14908 11812
rect 14973 11752 14986 11812
rect 14913 11711 14975 11719
rect 15020 11711 15027 11765
rect 15079 11711 15086 11765
rect 14913 11677 14926 11711
rect 14960 11682 14975 11711
rect 17044 11698 17096 11704
rect 14960 11677 17044 11682
rect 14913 11654 17044 11677
rect 17044 11631 17096 11637
rect 14531 11533 14540 11595
rect 14592 11533 14598 11595
rect 14934 11483 15143 11484
rect 14930 11468 15143 11483
rect 17255 11483 17308 11489
rect 14930 11456 17255 11468
rect 14930 11440 14993 11456
rect 15115 11440 17255 11456
rect 14930 11381 14962 11440
rect 14915 11374 14973 11381
rect 15021 11374 15027 11428
rect 15080 11374 15087 11428
rect 17255 11418 17308 11424
rect 14915 11340 14927 11374
rect 14961 11340 14973 11374
rect 14915 11330 14973 11340
rect 14533 11196 14540 11256
rect 14592 11196 14599 11256
rect 14903 11240 14915 11298
rect 14976 11240 14988 11298
<< via1 >>
rect 16975 13051 17027 13103
rect 17185 12671 17237 12728
rect 15008 12421 15060 12473
rect 17115 12415 17167 12474
rect 14533 12035 14595 12103
rect 16906 12039 16958 12093
rect 14908 11800 14973 11812
rect 14908 11764 14926 11800
rect 14926 11764 14961 11800
rect 14961 11764 14973 11800
rect 14908 11752 14973 11764
rect 15027 11755 15079 11765
rect 15027 11721 15036 11755
rect 15036 11721 15070 11755
rect 15070 11721 15079 11755
rect 15027 11711 15079 11721
rect 17044 11637 17096 11698
rect 14540 11579 14592 11595
rect 14540 11543 14547 11579
rect 14547 11543 14583 11579
rect 14583 11543 14592 11579
rect 14540 11533 14592 11543
rect 15027 11418 15080 11428
rect 15027 11384 15037 11418
rect 15037 11384 15071 11418
rect 15071 11384 15080 11418
rect 15027 11374 15080 11384
rect 17255 11424 17308 11483
rect 14540 11240 14592 11256
rect 14540 11206 14549 11240
rect 14549 11206 14583 11240
rect 14583 11206 14592 11240
rect 14540 11196 14592 11206
rect 14915 11286 14976 11298
rect 14915 11252 14927 11286
rect 14927 11252 14961 11286
rect 14961 11252 14976 11286
rect 14915 11240 14976 11252
<< metal2 >>
rect 15002 12421 15008 12473
rect 15060 12421 15066 12473
rect 14533 12103 14595 12110
rect 14533 12028 14595 12035
rect 14548 11595 14582 12028
rect 14900 11752 14908 11812
rect 14973 11752 14986 11812
rect 15020 11765 15063 12421
rect 14531 11533 14540 11595
rect 14592 11533 14598 11595
rect 14549 11256 14582 11533
rect 14926 11298 14964 11752
rect 15020 11711 15027 11765
rect 15079 11711 15086 11765
rect 15037 11428 15070 11711
rect 15021 11374 15027 11428
rect 15080 11374 15087 11428
rect 14533 11196 14540 11256
rect 14592 11196 14599 11256
rect 14903 11240 14915 11298
rect 14976 11240 14988 11298
rect 16846 9072 16876 15110
rect 16916 12099 16946 15115
rect 16986 13109 17016 15115
rect 16975 13103 17027 13109
rect 16975 13045 17027 13051
rect 16906 12093 16958 12099
rect 16906 12033 16958 12039
rect 16916 9077 16946 12033
rect 16986 9077 17016 13045
rect 17056 11704 17086 15114
rect 17126 12480 17156 15113
rect 17196 12734 17226 15109
rect 17185 12728 17237 12734
rect 17185 12665 17237 12671
rect 17115 12474 17167 12480
rect 17115 12409 17167 12415
rect 17044 11698 17096 11704
rect 17044 11631 17096 11637
rect 17056 9076 17086 11631
rect 17126 9075 17156 12409
rect 17196 9071 17226 12665
rect 17266 11489 17296 15114
rect 17255 11483 17308 11489
rect 17255 11418 17308 11424
rect 17266 9076 17296 11418
use lo_gen  lo_gen_0
timestamp 1647910564
transform 1 0 1884 0 1 7382
box 0 1500 10882 7765
use clk_tree  clk_tree_0 ~/cochlea_latest/fossi_cochlea/mag/clkgen
timestamp 1647885779
transform 0 1 -14948 -1 0 22337
box 0 0 18561 6322
use filter_p_m_fin  filter_p_m_fin_1
timestamp 1647909829
transform 1 0 5620 0 -1 21476
box -5284 -10468 28186 6398
use filter_p_m_fin  filter_p_m_fin_0
timestamp 1647909829
transform 1 0 5620 0 1 2680
box -5284 -10468 28186 6398
use filter_clkgen  filter_clkgen_0 ~/cochlea_latest/fossi_cochlea/mag/clkgen
timestamp 1647878126
transform 1 0 15039 0 1 11191
box -1895 666 1540 2096
use mux  mux_0
timestamp 1647510647
transform 0 -1 14944 1 0 11637
box -118 -152 220 422
use mux  mux_1
timestamp 1647510647
transform 0 -1 14945 1 0 11300
box -118 -152 220 422
<< labels >>
rlabel metal2 17283 9078 17283 9078 1 thresh_m
rlabel metal2 17071 9078 17071 9078 3 thresh_p
rlabel metal2 16862 9078 16862 9078 1 VDD
rlabel metal2 16930 9078 16930 9078 1 phi1
rlabel metal2 17001 9078 17001 9078 1 phi2
rlabel metal2 17139 9078 17139 9078 1 phi1b
rlabel metal2 17211 9078 17211 9078 1 phi2b
rlabel metal1 16579 13078 16579 13078 3 phi2
rlabel metal1 16557 12699 16557 12699 3 phi2b
rlabel metal1 16557 12447 16557 12447 3 phi1b
rlabel metal1 16579 12066 16579 12066 3 phi1
<< end >>
