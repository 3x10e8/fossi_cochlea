magic
tech sky130B
magscale 1 2
timestamp 1662788825
<< obsli1 >>
rect 1104 2159 94852 17425
<< obsm1 >>
rect 1104 2128 95206 17536
<< metal2 >>
rect 4434 19200 4490 20000
rect 12346 19200 12402 20000
rect 20258 19200 20314 20000
rect 28170 19200 28226 20000
rect 36082 19200 36138 20000
rect 43994 19200 44050 20000
rect 51906 19200 51962 20000
rect 59818 19200 59874 20000
rect 67730 19200 67786 20000
rect 75642 19200 75698 20000
rect 83554 19200 83610 20000
rect 91466 19200 91522 20000
rect 4434 0 4490 800
rect 12346 0 12402 800
rect 20258 0 20314 800
rect 28170 0 28226 800
rect 36082 0 36138 800
rect 43994 0 44050 800
rect 51906 0 51962 800
rect 59818 0 59874 800
rect 67730 0 67786 800
rect 75642 0 75698 800
rect 83554 0 83610 800
rect 91466 0 91522 800
<< obsm2 >>
rect 1582 19144 4378 19200
rect 4546 19144 12290 19200
rect 12458 19144 20202 19200
rect 20370 19144 28114 19200
rect 28282 19144 36026 19200
rect 36194 19144 43938 19200
rect 44106 19144 51850 19200
rect 52018 19144 59762 19200
rect 59930 19144 67674 19200
rect 67842 19144 75586 19200
rect 75754 19144 83498 19200
rect 83666 19144 91410 19200
rect 91578 19144 95202 19200
rect 1582 856 95202 19144
rect 1582 800 4378 856
rect 4546 800 12290 856
rect 12458 800 20202 856
rect 20370 800 28114 856
rect 28282 800 36026 856
rect 36194 800 43938 856
rect 44106 800 51850 856
rect 52018 800 59762 856
rect 59930 800 67674 856
rect 67842 800 75586 856
rect 75754 800 83498 856
rect 83666 800 91410 856
rect 91578 800 95202 856
<< metal3 >>
rect 95200 17280 96000 17400
rect 0 16600 800 16720
rect 95200 12384 96000 12504
rect 0 9936 800 10056
rect 95200 7488 96000 7608
rect 0 3272 800 3392
rect 95200 2592 96000 2712
<< obsm3 >>
rect 800 17200 95120 17441
rect 800 16800 95434 17200
rect 880 16520 95434 16800
rect 800 12584 95434 16520
rect 800 12304 95120 12584
rect 800 10136 95434 12304
rect 880 9856 95434 10136
rect 800 7688 95434 9856
rect 800 7408 95120 7688
rect 800 3472 95434 7408
rect 880 3192 95434 3472
rect 800 2792 95434 3192
rect 800 2512 95120 2792
rect 800 2143 95434 2512
<< metal4 >>
rect 12662 2128 12982 17456
rect 24380 2128 24700 17456
rect 36099 2128 36419 17456
rect 47817 2128 48137 17456
rect 59536 2128 59856 17456
rect 71254 2128 71574 17456
rect 82973 2128 83293 17456
rect 94691 2128 95011 17456
<< obsm4 >>
rect 59307 4795 59456 13157
rect 59936 4795 63605 13157
<< labels >>
rlabel metal2 s 28170 19200 28226 20000 6 cclk_I[0]
port 1 nsew signal output
rlabel metal2 s 75642 19200 75698 20000 6 cclk_I[1]
port 2 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 clk_master
port 5 nsew signal input
rlabel metal2 s 20258 19200 20314 20000 6 clkdiv2_I[0]
port 6 nsew signal output
rlabel metal2 s 67730 19200 67786 20000 6 clkdiv2_I[1]
port 7 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 clkdiv2_Q[0]
port 8 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 clkdiv2_Q[1]
port 9 nsew signal output
rlabel metal2 s 43994 19200 44050 20000 6 comp_high_I[0]
port 10 nsew signal input
rlabel metal2 s 91466 19200 91522 20000 6 comp_high_I[1]
port 11 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 comp_high_Q[0]
port 12 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 comp_high_Q[1]
port 13 nsew signal input
rlabel metal2 s 4434 19200 4490 20000 6 cos_out[0]
port 14 nsew signal output
rlabel metal2 s 51906 19200 51962 20000 6 cos_out[1]
port 15 nsew signal output
rlabel metal2 s 12346 19200 12402 20000 6 fb1_I[0]
port 16 nsew signal output
rlabel metal2 s 59818 19200 59874 20000 6 fb1_I[1]
port 17 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 fb1_Q[0]
port 18 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 fb1_Q[1]
port 19 nsew signal output
rlabel metal2 s 36082 19200 36138 20000 6 phi1b_dig_I[0]
port 20 nsew signal input
rlabel metal2 s 83554 19200 83610 20000 6 phi1b_dig_I[1]
port 21 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 phi1b_dig_Q[0]
port 22 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 phi1b_dig_Q[1]
port 23 nsew signal input
rlabel metal3 s 95200 17280 96000 17400 6 read_out_I[0]
port 24 nsew signal output
rlabel metal3 s 95200 12384 96000 12504 6 read_out_I[1]
port 25 nsew signal output
rlabel metal3 s 95200 7488 96000 7608 6 read_out_Q[0]
port 26 nsew signal output
rlabel metal3 s 95200 2592 96000 2712 6 read_out_Q[1]
port 27 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 rstb
port 28 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 sin_out[0]
port 29 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 sin_out[1]
port 30 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 ud_en
port 31 nsew signal input
rlabel metal4 s 12662 2128 12982 17456 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 36099 2128 36419 17456 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 59536 2128 59856 17456 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 82973 2128 83293 17456 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 24380 2128 24700 17456 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 47817 2128 48137 17456 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 71254 2128 71574 17456 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 94691 2128 95011 17456 6 vssd1
port 33 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 96000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4093632
string GDS_FILE /local_disk/fossi_cochlea/openlane/digital_unison/runs/22_09_09_22_44/results/signoff/digital_unison.magic.gds
string GDS_START 501876
<< end >>

