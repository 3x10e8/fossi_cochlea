magic
tech sky130A
magscale 1 2
timestamp 1654752206
<< obsli1 >>
rect 1104 2159 96876 77809
<< obsm1 >>
rect 1104 2128 96876 77840
<< metal2 >>
rect 2594 79200 2650 80000
rect 7746 79200 7802 80000
rect 12898 79200 12954 80000
rect 18050 79200 18106 80000
rect 23202 79200 23258 80000
rect 28354 79200 28410 80000
rect 33506 79200 33562 80000
rect 38658 79200 38714 80000
rect 43810 79200 43866 80000
rect 48962 79200 49018 80000
rect 54114 79200 54170 80000
rect 59266 79200 59322 80000
rect 64418 79200 64474 80000
rect 69570 79200 69626 80000
rect 74722 79200 74778 80000
rect 79874 79200 79930 80000
rect 85026 79200 85082 80000
rect 90178 79200 90234 80000
rect 95330 79200 95386 80000
rect 2686 0 2742 800
rect 8114 0 8170 800
rect 13542 0 13598 800
rect 18970 0 19026 800
rect 24398 0 24454 800
rect 29826 0 29882 800
rect 35346 0 35402 800
rect 40774 0 40830 800
rect 46202 0 46258 800
rect 51630 0 51686 800
rect 57058 0 57114 800
rect 62486 0 62542 800
rect 68006 0 68062 800
rect 73434 0 73490 800
rect 78862 0 78918 800
rect 84290 0 84346 800
rect 89718 0 89774 800
rect 95146 0 95202 800
<< obsm2 >>
rect 1398 79144 2538 79200
rect 2706 79144 7690 79200
rect 7858 79144 12842 79200
rect 13010 79144 17994 79200
rect 18162 79144 23146 79200
rect 23314 79144 28298 79200
rect 28466 79144 33450 79200
rect 33618 79144 38602 79200
rect 38770 79144 43754 79200
rect 43922 79144 48906 79200
rect 49074 79144 54058 79200
rect 54226 79144 59210 79200
rect 59378 79144 64362 79200
rect 64530 79144 69514 79200
rect 69682 79144 74666 79200
rect 74834 79144 79818 79200
rect 79986 79144 84970 79200
rect 85138 79144 90122 79200
rect 90290 79144 95274 79200
rect 95442 79144 96682 79200
rect 1398 856 96682 79144
rect 1398 734 2630 856
rect 2798 734 8058 856
rect 8226 734 13486 856
rect 13654 734 18914 856
rect 19082 734 24342 856
rect 24510 734 29770 856
rect 29938 734 35290 856
rect 35458 734 40718 856
rect 40886 734 46146 856
rect 46314 734 51574 856
rect 51742 734 57002 856
rect 57170 734 62430 856
rect 62598 734 67950 856
rect 68118 734 73378 856
rect 73546 734 78806 856
rect 78974 734 84234 856
rect 84402 734 89662 856
rect 89830 734 95090 856
rect 95258 734 96682 856
<< metal3 >>
rect 0 77664 800 77784
rect 97200 77800 98000 77920
rect 97200 73584 98000 73704
rect 0 73176 800 73296
rect 97200 69368 98000 69488
rect 0 68824 800 68944
rect 97200 65152 98000 65272
rect 0 64336 800 64456
rect 97200 60936 98000 61056
rect 0 59848 800 59968
rect 97200 56720 98000 56840
rect 0 55496 800 55616
rect 97200 52504 98000 52624
rect 0 51008 800 51128
rect 97200 48288 98000 48408
rect 0 46520 800 46640
rect 97200 44072 98000 44192
rect 0 42168 800 42288
rect 97200 39856 98000 39976
rect 0 37680 800 37800
rect 97200 35640 98000 35760
rect 0 33192 800 33312
rect 97200 31424 98000 31544
rect 0 28840 800 28960
rect 97200 27208 98000 27328
rect 0 24352 800 24472
rect 97200 22992 98000 23112
rect 0 19864 800 19984
rect 97200 18776 98000 18896
rect 0 15512 800 15632
rect 97200 14560 98000 14680
rect 0 11024 800 11144
rect 97200 10344 98000 10464
rect 0 6536 800 6656
rect 97200 6128 98000 6248
rect 0 2184 800 2304
rect 97200 2048 98000 2168
<< obsm3 >>
rect 800 77864 97120 77890
rect 880 77720 97120 77864
rect 880 77584 97200 77720
rect 800 73784 97200 77584
rect 800 73504 97120 73784
rect 800 73376 97200 73504
rect 880 73096 97200 73376
rect 800 69568 97200 73096
rect 800 69288 97120 69568
rect 800 69024 97200 69288
rect 880 68744 97200 69024
rect 800 65352 97200 68744
rect 800 65072 97120 65352
rect 800 64536 97200 65072
rect 880 64256 97200 64536
rect 800 61136 97200 64256
rect 800 60856 97120 61136
rect 800 60048 97200 60856
rect 880 59768 97200 60048
rect 800 56920 97200 59768
rect 800 56640 97120 56920
rect 800 55696 97200 56640
rect 880 55416 97200 55696
rect 800 52704 97200 55416
rect 800 52424 97120 52704
rect 800 51208 97200 52424
rect 880 50928 97200 51208
rect 800 48488 97200 50928
rect 800 48208 97120 48488
rect 800 46720 97200 48208
rect 880 46440 97200 46720
rect 800 44272 97200 46440
rect 800 43992 97120 44272
rect 800 42368 97200 43992
rect 880 42088 97200 42368
rect 800 40056 97200 42088
rect 800 39776 97120 40056
rect 800 37880 97200 39776
rect 880 37600 97200 37880
rect 800 35840 97200 37600
rect 800 35560 97120 35840
rect 800 33392 97200 35560
rect 880 33112 97200 33392
rect 800 31624 97200 33112
rect 800 31344 97120 31624
rect 800 29040 97200 31344
rect 880 28760 97200 29040
rect 800 27408 97200 28760
rect 800 27128 97120 27408
rect 800 24552 97200 27128
rect 880 24272 97200 24552
rect 800 23192 97200 24272
rect 800 22912 97120 23192
rect 800 20064 97200 22912
rect 880 19784 97200 20064
rect 800 18976 97200 19784
rect 800 18696 97120 18976
rect 800 15712 97200 18696
rect 880 15432 97200 15712
rect 800 14760 97200 15432
rect 800 14480 97120 14760
rect 800 11224 97200 14480
rect 880 10944 97200 11224
rect 800 10544 97200 10944
rect 800 10264 97120 10544
rect 800 6736 97200 10264
rect 880 6456 97200 6736
rect 800 6328 97200 6456
rect 800 6048 97120 6328
rect 800 2384 97200 6048
rect 880 2248 97200 2384
rect 880 2104 97120 2248
rect 800 2075 97120 2104
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
rect 81008 2128 81328 77840
rect 96368 2128 96688 77840
<< obsm4 >>
rect 20483 2347 34848 72589
rect 35328 2347 50208 72589
rect 50688 2347 65568 72589
rect 66048 2347 80928 72589
rect 81408 2347 89733 72589
<< labels >>
rlabel metal3 s 0 24352 800 24472 6 cclk_I[0]
port 1 nsew signal output
rlabel metal3 s 0 55496 800 55616 6 cclk_I[1]
port 2 nsew signal output
rlabel metal3 s 97200 6128 98000 6248 6 cclk_Q[0]
port 3 nsew signal output
rlabel metal3 s 97200 35640 98000 35760 6 cclk_Q[1]
port 4 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 clk_master
port 5 nsew signal input
rlabel metal2 s 7746 79200 7802 80000 6 clk_master_out
port 6 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 clkdiv2_I[0]
port 7 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 clkdiv2_I[1]
port 8 nsew signal output
rlabel metal3 s 97200 10344 98000 10464 6 clkdiv2_Q[0]
port 9 nsew signal output
rlabel metal3 s 97200 39856 98000 39976 6 clkdiv2_Q[1]
port 10 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 clkdiv2_in
port 11 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 comp_high_I[0]
port 12 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 comp_high_I[1]
port 13 nsew signal input
rlabel metal3 s 97200 14560 98000 14680 6 comp_high_Q[0]
port 14 nsew signal input
rlabel metal3 s 97200 44072 98000 44192 6 comp_high_Q[1]
port 15 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 cos_out[0]
port 16 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 cos_out[1]
port 17 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 cos_outb[0]
port 18 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 cos_outb[1]
port 19 nsew signal output
rlabel metal2 s 18050 79200 18106 80000 6 div2out
port 20 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 fb1_I[0]
port 21 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 fb1_I[1]
port 22 nsew signal output
rlabel metal3 s 97200 22992 98000 23112 6 fb1_Q[0]
port 23 nsew signal output
rlabel metal3 s 97200 52504 98000 52624 6 fb1_Q[1]
port 24 nsew signal output
rlabel metal3 s 97200 69368 98000 69488 6 fb2_I[0]
port 25 nsew signal output
rlabel metal3 s 97200 73584 98000 73704 6 fb2_I[1]
port 26 nsew signal output
rlabel metal3 s 0 73176 800 73296 6 fb2_Q[0]
port 27 nsew signal output
rlabel metal3 s 97200 77800 98000 77920 6 fb2_Q[1]
port 28 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 gray_clk_in[0]
port 29 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 gray_clk_in[1]
port 30 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 gray_clk_in[2]
port 31 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 gray_clk_in[3]
port 32 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 gray_clk_in[4]
port 33 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 gray_clk_in[5]
port 34 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 gray_clk_in[6]
port 35 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 gray_clk_in[7]
port 36 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 gray_clk_in[8]
port 37 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 gray_clk_in[9]
port 38 nsew signal input
rlabel metal2 s 69570 79200 69626 80000 6 gray_clk_out[10]
port 39 nsew signal output
rlabel metal2 s 23202 79200 23258 80000 6 gray_clk_out[1]
port 40 nsew signal output
rlabel metal2 s 28354 79200 28410 80000 6 gray_clk_out[2]
port 41 nsew signal output
rlabel metal2 s 33506 79200 33562 80000 6 gray_clk_out[3]
port 42 nsew signal output
rlabel metal2 s 38658 79200 38714 80000 6 gray_clk_out[4]
port 43 nsew signal output
rlabel metal2 s 43810 79200 43866 80000 6 gray_clk_out[5]
port 44 nsew signal output
rlabel metal2 s 48962 79200 49018 80000 6 gray_clk_out[6]
port 45 nsew signal output
rlabel metal2 s 54114 79200 54170 80000 6 gray_clk_out[7]
port 46 nsew signal output
rlabel metal2 s 59266 79200 59322 80000 6 gray_clk_out[8]
port 47 nsew signal output
rlabel metal2 s 64418 79200 64474 80000 6 gray_clk_out[9]
port 48 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 no_ones_below_in[0]
port 49 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 no_ones_below_in[1]
port 50 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 no_ones_below_in[2]
port 51 nsew signal input
rlabel metal2 s 74722 79200 74778 80000 6 no_ones_below_out[0]
port 52 nsew signal output
rlabel metal2 s 79874 79200 79930 80000 6 no_ones_below_out[1]
port 53 nsew signal output
rlabel metal2 s 85026 79200 85082 80000 6 no_ones_below_out[2]
port 54 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 phi1b_dig_I[0]
port 55 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 phi1b_dig_I[1]
port 56 nsew signal input
rlabel metal3 s 97200 18776 98000 18896 6 phi1b_dig_Q[0]
port 57 nsew signal input
rlabel metal3 s 97200 48288 98000 48408 6 phi1b_dig_Q[1]
port 58 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 read_out_I[0]
port 59 nsew signal output
rlabel metal2 s 95330 79200 95386 80000 6 read_out_I[1]
port 60 nsew signal output
rlabel metal3 s 0 64336 800 64456 6 read_out_I_top[0]
port 61 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 read_out_I_top[1]
port 62 nsew signal output
rlabel metal2 s 90178 79200 90234 80000 6 read_out_Q[0]
port 63 nsew signal output
rlabel metal3 s 0 77664 800 77784 6 read_out_Q[1]
port 64 nsew signal output
rlabel metal3 s 97200 60936 98000 61056 6 read_out_Q_top[0]
port 65 nsew signal output
rlabel metal3 s 97200 65152 98000 65272 6 read_out_Q_top[1]
port 66 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 rstb
port 67 nsew signal input
rlabel metal2 s 2594 79200 2650 80000 6 rstb_out
port 68 nsew signal output
rlabel metal3 s 97200 2048 98000 2168 6 sin_out[0]
port 69 nsew signal output
rlabel metal3 s 97200 31424 98000 31544 6 sin_out[1]
port 70 nsew signal output
rlabel metal3 s 97200 27208 98000 27328 6 sin_outb[0]
port 71 nsew signal output
rlabel metal3 s 97200 56720 98000 56840 6 sin_outb[1]
port 72 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 ud_en
port 73 nsew signal input
rlabel metal2 s 12898 79200 12954 80000 6 ud_en_out
port 74 nsew signal output
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 75 nsew power input
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 75 nsew power input
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 75 nsew power input
rlabel metal4 s 96368 2128 96688 77840 6 vccd1
port 75 nsew power input
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 76 nsew ground input
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 76 nsew ground input
rlabel metal4 s 81008 2128 81328 77840 6 vssd1
port 76 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 98000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8201018
string GDS_FILE /Volumes/export/isn/abhinav/fossi_cochlea/openlane/scalable_dual_core/runs/scalable_dual_core/results/finishing/scalable_dual_core.magic.gds
string GDS_START 415174
<< end >>

