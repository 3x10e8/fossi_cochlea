magic
tech sky130B
magscale 1 2
timestamp 1663892726
<< nwell >>
rect 25556 34014 25620 34078
<< psubdiff >>
rect 25260 33477 25311 33527
<< locali >>
rect 25260 33477 25311 33527
rect 22218 28813 22252 29386
rect 25824 28777 25858 29363
<< viali >>
rect 22218 29386 22252 29420
<< metal1 >>
rect 18870 35470 18934 35476
rect 18870 35418 18876 35470
rect 18928 35461 18934 35470
rect 21976 35461 21982 35470
rect 18928 35427 21982 35461
rect 18928 35418 18934 35427
rect 21976 35418 21982 35427
rect 22034 35418 22040 35470
rect 18870 35412 18934 35418
rect 5046 35088 5052 35140
rect 5104 35131 5110 35140
rect 8874 35131 8880 35140
rect 5104 35097 8880 35131
rect 5104 35088 5110 35097
rect 8874 35088 8880 35097
rect 8932 35088 8938 35140
rect 24646 34878 24698 34884
rect 23265 34828 24646 34872
rect 24646 34820 24698 34826
rect 8490 34372 8768 34468
rect 9858 34464 11514 34468
rect 9858 34376 11276 34464
rect 11508 34376 11514 34464
rect 36790 34464 38446 34468
rect 24403 34390 24455 34396
rect 9858 34372 11514 34376
rect 8490 33380 8590 34372
rect 23252 34341 24403 34385
rect 36790 34376 36796 34464
rect 37028 34376 38446 34464
rect 36790 34372 38446 34376
rect 39536 34372 39814 34468
rect 24403 34332 24455 34338
rect 23531 34021 24319 34100
rect 25556 34071 25620 34078
rect 25556 34019 25562 34071
rect 25614 34019 25620 34071
rect 25556 34014 25620 34019
rect 8642 33924 8812 33930
rect 39492 33924 39662 33930
rect 19238 33892 19270 33900
rect 8642 33822 8812 33828
rect 19130 33810 19270 33892
rect 39492 33822 39662 33828
rect 19238 33474 19270 33810
rect 24210 33769 24262 33775
rect 23256 33721 24210 33765
rect 24210 33711 24262 33717
rect 22302 33656 22308 33665
rect 22099 33622 22308 33656
rect 22302 33613 22308 33622
rect 22360 33613 22366 33665
rect 23547 33479 24335 33558
rect 25260 33477 25311 33527
rect 39714 33380 39814 34372
rect 8490 33284 8798 33380
rect 23757 33297 23810 33303
rect 23250 33253 23757 33297
rect 26380 33297 26456 33303
rect 23810 33245 24300 33291
rect 23757 33239 24300 33245
rect 23789 33237 24300 33239
rect 26380 33233 26386 33297
rect 26450 33233 26456 33297
rect 39506 33284 39814 33380
rect 26380 33227 26456 33233
rect 13512 32980 13518 33032
rect 13570 33023 13576 33032
rect 13570 33022 13746 33023
rect 13570 32989 18702 33022
rect 13570 32980 13576 32989
rect 13746 32988 18702 32989
rect 23538 32927 24326 33006
rect 23593 32672 23646 32678
rect 23229 32615 23593 32672
rect 23645 32615 23646 32672
rect 23593 32609 23646 32615
rect 23225 32270 23277 32276
rect 23225 32103 23277 32109
rect 38286 30304 38292 30356
rect 38344 30304 38350 30356
rect 37773 30236 37825 30242
rect 37773 30178 37825 30184
rect 24402 30120 24456 30126
rect 24402 30068 24403 30120
rect 24455 30068 24456 30120
rect 24402 30062 24456 30068
rect 24645 29997 24697 30003
rect 24645 29939 24697 29945
rect 23758 29880 23810 29886
rect 23758 29822 23810 29828
rect 24209 29756 24261 29762
rect 24209 29698 24261 29704
rect 23593 28713 23645 28719
rect 22201 28666 23593 28711
rect 23645 28666 25876 28711
rect 23593 28654 23645 28661
rect 23224 28544 23276 28550
rect 22279 28496 23224 28541
rect 23276 28496 25793 28541
rect 23224 28486 23276 28492
rect 24645 28453 24697 28459
rect 23390 28447 23442 28453
rect 22206 28406 23390 28440
rect 23442 28406 24645 28440
rect 24697 28406 25871 28440
rect 24645 28395 24697 28401
rect 23390 28389 23442 28395
rect 23878 27615 23884 27624
rect 22284 27581 23884 27615
rect 22284 26349 22318 27581
rect 23878 27572 23884 27581
rect 23936 27572 23942 27624
<< via1 >>
rect 18876 35418 18928 35470
rect 21982 35418 22034 35470
rect 5052 35088 5104 35140
rect 8880 35088 8932 35140
rect 24646 34826 24698 34878
rect 11276 34376 11508 34464
rect 24403 34338 24455 34390
rect 36796 34376 37028 34464
rect 25562 34019 25614 34071
rect 8642 33828 8812 33924
rect 39492 33828 39662 33924
rect 24210 33717 24262 33769
rect 26207 33714 26259 33766
rect 22308 33613 22360 33665
rect 8962 33292 9194 33370
rect 10676 33292 10908 33370
rect 23757 33245 23810 33297
rect 26386 33233 26450 33297
rect 37396 33292 37628 33370
rect 39110 33292 39342 33370
rect 13518 32980 13570 33032
rect 25478 32918 25690 33006
rect 23593 32615 23645 32672
rect 23225 32109 23277 32270
rect 38292 30304 38344 30356
rect 37773 30184 37825 30236
rect 24403 30068 24455 30120
rect 24645 29945 24697 29997
rect 23758 29828 23810 29880
rect 24209 29704 24261 29756
rect 23593 28661 23645 28713
rect 23224 28492 23276 28544
rect 23390 28395 23442 28447
rect 24645 28401 24697 28453
rect 23884 27572 23936 27624
rect 24018 26706 24070 26758
<< metal2 >>
rect 5052 35140 5108 37140
rect 5104 35088 5108 35140
rect 5052 35082 5108 35088
rect 8880 35140 8932 35146
rect 8880 35082 8932 35088
rect 8642 33924 8812 33930
rect 8642 29658 8812 33828
rect 8889 33650 8923 35082
rect 11276 34464 11508 34470
rect 8962 33370 9194 33380
rect 8962 30998 9194 33292
rect 9969 31160 10003 33860
rect 10488 31336 10522 33848
rect 10676 33370 10908 33380
rect 10460 31328 10550 31336
rect 10460 31258 10470 31328
rect 10540 31258 10550 31328
rect 10460 31250 10550 31258
rect 9940 31152 10030 31160
rect 9940 31082 9950 31152
rect 10020 31082 10030 31152
rect 9940 31074 10030 31082
rect 8952 30990 9204 30998
rect 8952 30886 8962 30990
rect 9194 30886 9204 30990
rect 8952 30876 9204 30886
rect 8600 29648 8852 29658
rect 10676 29656 10908 33292
rect 8600 29550 8610 29648
rect 8842 29550 8852 29648
rect 8600 29540 8852 29550
rect 10666 29648 10918 29656
rect 10666 29550 10676 29648
rect 10908 29550 10918 29648
rect 10666 29540 10918 29550
rect 11276 29472 11508 34376
rect 13516 33032 13572 37140
rect 18870 35470 18934 35476
rect 18870 35418 18876 35470
rect 18928 35418 18934 35470
rect 18870 35412 18934 35418
rect 21980 35470 22036 37140
rect 30444 35490 30500 37140
rect 21980 35418 21982 35470
rect 22034 35418 22036 35470
rect 21980 35416 22036 35418
rect 30429 35481 30511 35490
rect 21982 35412 22034 35416
rect 18885 33952 18919 35412
rect 30429 35409 30434 35481
rect 30506 35409 30511 35481
rect 30429 35404 30511 35409
rect 33938 35459 34002 35468
rect 38908 35466 38964 37140
rect 30434 35400 30506 35404
rect 24646 34878 24698 34884
rect 24646 34820 24698 34826
rect 24403 34390 24455 34396
rect 13516 32980 13518 33032
rect 13570 32980 13572 33032
rect 13516 32979 13572 32980
rect 13518 32974 13570 32979
rect 21478 31727 21508 34350
rect 24403 34332 24455 34338
rect 24210 33769 24262 33775
rect 24210 33711 24262 33717
rect 22308 33665 22360 33671
rect 22308 33607 22360 33613
rect 21463 31718 21523 31727
rect 21463 31649 21523 31658
rect 22317 31523 22351 33607
rect 23757 33297 23810 33303
rect 23757 33239 23810 33245
rect 23593 32672 23646 32678
rect 23645 32615 23646 32672
rect 23593 32609 23646 32615
rect 23225 32270 23277 32276
rect 23225 32103 23277 32109
rect 22304 31514 22364 31523
rect 22304 31445 22364 31454
rect 21701 30758 21757 30767
rect 21701 30693 21757 30702
rect 21714 30481 21748 30693
rect 22096 30579 22130 30580
rect 22085 30570 22141 30579
rect 22085 30505 22141 30514
rect 11266 29456 11518 29472
rect 11266 29358 11276 29456
rect 11508 29358 11518 29456
rect 11266 29348 11518 29358
rect 21713 28443 21749 30481
rect 21713 28405 21922 28443
rect 22095 28442 22131 30505
rect 22202 28666 22240 28717
rect 23227 28551 23275 32103
rect 23594 28719 23644 32609
rect 23758 29880 23810 33239
rect 23758 29809 23810 29828
rect 24009 30958 24080 30970
rect 24009 30902 24017 30958
rect 24073 30902 24080 30958
rect 23593 28713 23645 28719
rect 23593 28654 23645 28661
rect 23224 28544 23276 28551
rect 23224 28486 23276 28492
rect 23390 28447 23442 28453
rect 23390 28389 23442 28395
rect 23400 26902 23434 28389
rect 23884 27624 23936 27630
rect 23865 27567 23874 27623
rect 23936 27572 23939 27623
rect 23930 27567 23939 27572
rect 23884 27566 23936 27567
rect 24009 26758 24080 30902
rect 24211 29762 24260 33711
rect 24404 30126 24454 34332
rect 24402 30120 24456 30126
rect 24402 30068 24403 30120
rect 24455 30068 24456 30120
rect 24402 30062 24456 30068
rect 24404 30060 24454 30062
rect 24647 30003 24696 34820
rect 25560 34075 25618 34084
rect 25560 34008 25618 34017
rect 26195 33774 26275 33783
rect 26195 33711 26204 33774
rect 26266 33711 26275 33774
rect 26195 33702 26275 33711
rect 26380 33297 26456 33303
rect 26380 33233 26386 33297
rect 26450 33233 26456 33297
rect 26380 33227 26456 33233
rect 25468 33006 25700 33014
rect 25468 32918 25478 33006
rect 25690 32918 25700 33006
rect 25468 30986 25700 32918
rect 26386 32115 26450 33227
rect 33938 32119 34002 35395
rect 38906 35457 38966 35466
rect 38906 35388 38966 35397
rect 39368 34985 39428 34994
rect 47372 34992 47428 37140
rect 47368 34983 47428 34992
rect 47368 34927 47370 34983
rect 47426 34927 47428 34983
rect 47368 34925 47428 34927
rect 39368 34916 39428 34925
rect 47370 34918 47426 34925
rect 36796 34464 37028 34470
rect 26386 32042 26450 32051
rect 33934 32113 34006 32119
rect 33934 32057 33942 32113
rect 33998 32057 34006 32113
rect 33934 32048 34006 32057
rect 25468 30886 25474 30986
rect 25694 30886 25700 30986
rect 25468 30876 25700 30886
rect 25935 30765 25991 30774
rect 25935 30700 25991 30709
rect 24645 29997 24697 30003
rect 24645 29939 24697 29945
rect 24647 29925 24696 29939
rect 24209 29756 24261 29762
rect 24209 29698 24261 29704
rect 25820 28683 25861 28717
rect 24645 28453 24697 28459
rect 25946 28432 25980 30700
rect 26315 30568 26371 30578
rect 26315 30503 26371 30512
rect 26328 28440 26362 30503
rect 36796 29472 37028 34376
rect 37396 33370 37628 33380
rect 37396 29656 37628 33292
rect 37782 30236 37816 33852
rect 38301 30362 38335 33864
rect 39381 33650 39415 34916
rect 39492 33924 39662 33930
rect 39110 33370 39342 33380
rect 39110 30998 39342 33292
rect 39100 30990 39352 30998
rect 39100 30886 39110 30990
rect 39342 30886 39352 30990
rect 39100 30876 39352 30886
rect 38292 30356 38344 30362
rect 38292 30298 38344 30304
rect 37767 30184 37773 30236
rect 37825 30184 37831 30236
rect 39492 29658 39662 33828
rect 37386 29648 37638 29656
rect 37386 29550 37396 29648
rect 37628 29550 37638 29648
rect 37386 29540 37638 29550
rect 39452 29648 39704 29658
rect 39452 29550 39462 29648
rect 39694 29550 39704 29648
rect 39452 29540 39704 29550
rect 36786 29456 37038 29472
rect 36786 29358 36796 29456
rect 37028 29358 37038 29456
rect 36786 29348 37038 29358
rect 26152 28403 26362 28440
rect 24645 28395 24697 28401
rect 24656 26902 24690 28395
rect 24009 26706 24018 26758
rect 24070 26706 24080 26758
rect 24009 26700 24080 26706
rect 46310 26270 47033 26314
rect 24015 26077 24071 26081
rect 46310 26064 46355 26270
rect 1063 26007 1751 26051
<< via2 >>
rect 10470 31258 10540 31328
rect 9950 31082 10020 31152
rect 8962 30886 9194 30990
rect 8610 29550 8842 29648
rect 10676 29550 10908 29648
rect 30434 35409 30506 35481
rect 33938 35395 34002 35459
rect 21463 31658 21523 31718
rect 22304 31454 22364 31514
rect 21701 30702 21757 30758
rect 22085 30514 22141 30570
rect 11276 29358 11508 29456
rect 24017 30902 24073 30958
rect 23874 27572 23884 27623
rect 23884 27572 23930 27623
rect 23874 27567 23930 27572
rect 25560 34071 25618 34075
rect 25560 34019 25562 34071
rect 25562 34019 25614 34071
rect 25614 34019 25618 34071
rect 25560 34017 25618 34019
rect 26204 33766 26266 33774
rect 26204 33714 26207 33766
rect 26207 33714 26259 33766
rect 26259 33714 26266 33766
rect 26204 33711 26266 33714
rect 25478 32918 25690 33006
rect 38906 35397 38966 35457
rect 39368 34925 39428 34985
rect 47370 34927 47426 34983
rect 26386 32051 26450 32115
rect 33942 32057 33998 32113
rect 25474 30886 25694 30986
rect 25935 30709 25991 30765
rect 26315 30512 26371 30568
rect 39110 30886 39342 30990
rect 37396 29550 37628 29648
rect 39462 29550 39694 29648
rect 36796 29358 37028 29456
<< metal3 >>
rect 23866 35485 30511 35486
rect 23861 35405 23867 35485
rect 23947 35481 30511 35485
rect 23947 35409 30434 35481
rect 30506 35409 30511 35481
rect 23947 35405 30511 35409
rect 23866 35404 30511 35405
rect 33933 35459 34007 35464
rect 38901 35459 38971 35462
rect 33933 35395 33938 35459
rect 34002 35457 38971 35459
rect 34002 35397 38906 35457
rect 38966 35397 38971 35457
rect 34002 35395 38971 35397
rect 33933 35390 34007 35395
rect 38901 35392 38971 35395
rect 39363 34985 39433 34990
rect 47365 34985 47431 34988
rect 39363 34925 39368 34985
rect 39428 34983 47431 34985
rect 39428 34927 47370 34983
rect 47426 34927 47431 34983
rect 39428 34925 47431 34927
rect 39363 34920 39433 34925
rect 47365 34922 47431 34925
rect 25540 34078 25640 34095
rect 25540 34014 25556 34078
rect 25620 34014 25640 34078
rect 25540 33996 25640 34014
rect 26179 33783 26288 33800
rect 26179 33702 26195 33783
rect 26275 33702 26288 33783
rect 26179 33692 26288 33702
rect 25468 33006 25700 33014
rect 25468 32918 25478 33006
rect 25690 32918 25700 33006
rect 25468 32910 25700 32918
rect 26381 32117 26455 32120
rect 33937 32117 34003 32118
rect 24731 32053 24737 32117
rect 24801 32115 34003 32117
rect 24801 32053 26386 32115
rect 26381 32051 26386 32053
rect 26450 32113 34003 32115
rect 26450 32057 33942 32113
rect 33998 32057 34003 32113
rect 26450 32053 34003 32057
rect 26450 32051 26455 32053
rect 33937 32052 34003 32053
rect 26381 32046 26455 32051
rect -26 31718 50758 31740
rect -26 31658 21463 31718
rect 21523 31658 50758 31718
rect -26 31640 50758 31658
rect -26 31514 50758 31540
rect -26 31454 22304 31514
rect 22364 31454 50758 31514
rect -26 31440 50758 31454
rect 10460 31328 10550 31336
rect 5834 31324 5920 31326
rect 5834 31260 5840 31324
rect 5914 31322 5920 31324
rect 10460 31322 10470 31328
rect 5914 31262 10470 31322
rect 5914 31260 5920 31262
rect 5834 31258 5920 31260
rect 10460 31258 10470 31262
rect 10540 31258 10550 31328
rect 10460 31250 10550 31258
rect 9940 31152 10030 31160
rect 9940 31082 9950 31152
rect 10020 31146 10030 31152
rect 42156 31148 42242 31150
rect 42156 31146 42162 31148
rect 10020 31086 42162 31146
rect 10020 31082 10030 31086
rect 42156 31084 42162 31086
rect 42236 31084 42242 31148
rect 42156 31082 42242 31084
rect 9940 31074 10030 31082
rect 8952 30990 9204 30998
rect 8952 30986 8962 30990
rect -26 30886 8962 30986
rect 9194 30986 9204 30990
rect 25468 30986 25700 30996
rect 39100 30990 39352 30998
rect 39100 30986 39110 30990
rect 9194 30971 25474 30986
rect 9194 30895 18624 30971
rect 18710 30958 25474 30971
rect 18710 30902 24017 30958
rect 24073 30902 25474 30958
rect 18710 30895 25474 30902
rect 9194 30886 25474 30895
rect 25694 30886 39110 30986
rect 39342 30986 39352 30990
rect 39342 30886 50758 30986
rect 8952 30876 9204 30886
rect 25468 30876 25700 30886
rect 39100 30876 39352 30886
rect -26 30765 50758 30786
rect -26 30758 25935 30765
rect -26 30702 21701 30758
rect 21757 30709 25935 30758
rect 25991 30709 50758 30765
rect 21757 30702 50758 30709
rect -26 30686 50758 30702
rect -26 30570 50758 30586
rect -26 30514 22085 30570
rect 22141 30568 50758 30570
rect 22141 30514 26315 30568
rect -26 30512 26315 30514
rect 26371 30512 50758 30568
rect -26 30486 50758 30512
rect 8600 29649 8852 29658
rect 10666 29649 10918 29656
rect 37386 29649 37638 29656
rect 39452 29649 39704 29658
rect -26 29648 23388 29649
rect -26 29550 8610 29648
rect 8842 29550 10676 29648
rect 10908 29636 23388 29648
rect 10908 29565 22940 29636
rect 23014 29565 23388 29636
rect 10908 29550 23388 29565
rect -26 29549 23388 29550
rect 36482 29648 39862 29649
rect 36482 29550 37396 29648
rect 37628 29550 39462 29648
rect 39694 29550 39862 29648
rect 36482 29549 39862 29550
rect 46890 29549 50758 29649
rect 8600 29540 8852 29549
rect 10666 29540 10918 29549
rect 37386 29540 37638 29549
rect 39452 29540 39704 29549
rect -26 29358 492 29458
rect 11266 29456 11518 29472
rect 11266 29358 11276 29456
rect 11508 29358 11518 29456
rect 28122 29358 33044 29458
rect 36786 29456 37038 29472
rect 36786 29358 36796 29456
rect 37028 29358 37038 29456
rect 47584 29358 50758 29458
rect 11266 29348 11518 29358
rect 36786 29348 37038 29358
rect 23854 27633 23954 27642
rect 23854 27560 23871 27633
rect 23944 27560 23954 27633
rect 23854 27544 23954 27560
rect 23278 26637 23355 26642
rect 23278 26571 23284 26637
rect 23349 26571 23355 26637
rect 23278 26566 23355 26571
rect 24730 26636 24807 26642
rect 24730 26572 24737 26636
rect 24801 26572 24807 26636
rect 24730 26566 24807 26572
rect 24004 26083 24081 26092
rect 24004 26019 24010 26083
rect 24074 26019 24081 26083
rect 24004 26013 24081 26019
<< via3 >>
rect 23867 35405 23947 35485
rect 25556 34075 25620 34078
rect 25556 34017 25560 34075
rect 25560 34017 25618 34075
rect 25618 34017 25620 34075
rect 25556 34014 25620 34017
rect 26195 33774 26275 33783
rect 26195 33711 26204 33774
rect 26204 33711 26266 33774
rect 26266 33711 26275 33774
rect 26195 33702 26275 33711
rect 25478 32918 25690 33006
rect 24737 32053 24801 32117
rect 5840 31260 5914 31324
rect 42162 31084 42236 31148
rect 18624 30895 18710 30971
rect 22940 29565 23014 29636
rect 22483 29373 22555 29445
rect 23871 27623 23944 27633
rect 23871 27567 23874 27623
rect 23874 27567 23930 27623
rect 23930 27567 23944 27623
rect 23871 27560 23944 27567
rect 23284 26571 23349 26637
rect 24737 26572 24801 26636
rect 24010 26019 24074 26083
<< metal4 >>
rect 23866 35485 23948 35486
rect 23866 35405 23867 35485
rect 23947 35405 23948 35485
rect 23866 32739 23948 35405
rect 25550 34078 25625 34079
rect 25550 34014 25556 34078
rect 25620 34014 25625 34078
rect 25550 33014 25625 34014
rect 26179 33783 26288 33800
rect 26179 33777 26195 33783
rect 26043 33704 26195 33777
rect 25468 33006 25700 33014
rect 25468 32918 25478 33006
rect 25690 32918 25700 33006
rect 25468 32910 25700 32918
rect 5834 31324 5920 31326
rect 5834 31260 5840 31324
rect 5914 31260 5920 31324
rect 5834 31258 5920 31260
rect 5840 25993 5914 31258
rect 18618 30971 18716 32261
rect 18618 30895 18624 30971
rect 18710 30895 18716 30971
rect 18618 30886 18716 30895
rect 22481 29445 22558 31932
rect 22933 29636 23019 31843
rect 22933 29565 22940 29636
rect 23014 29565 23019 29636
rect 22933 29532 23019 29565
rect 22481 29373 22483 29445
rect 22555 29373 22558 29445
rect 22481 29341 22558 29373
rect 23870 27633 23945 32739
rect 26044 32504 26111 33704
rect 26179 33702 26195 33704
rect 26275 33702 26288 33783
rect 26179 33692 26288 33702
rect 23870 27560 23871 27633
rect 23944 27560 23945 27633
rect 23870 27559 23945 27560
rect 24241 32432 26111 32504
rect 24241 27210 24316 32432
rect 24736 32117 24802 32118
rect 24736 32053 24737 32117
rect 24801 32053 24802 32117
rect 24736 32052 24802 32053
rect 23824 27124 24316 27210
rect 23284 26642 23349 26769
rect 23278 26637 23355 26642
rect 23278 26571 23284 26637
rect 23349 26571 23355 26637
rect 23278 26566 23355 26571
rect 24010 26089 24076 27124
rect 24737 26642 24801 32052
rect 42156 31148 42242 31150
rect 42156 31084 42162 31148
rect 42236 31084 42242 31148
rect 42156 31082 42242 31084
rect 24730 26636 24807 26642
rect 24730 26572 24737 26636
rect 24801 26572 24807 26636
rect 24730 26566 24807 26572
rect 24004 26083 24081 26089
rect 24004 26019 24010 26083
rect 24074 26019 24081 26083
rect 24004 26013 24081 26019
rect 42162 25993 42236 31082
rect -26 961 1074 1160
rect 47129 961 50758 1160
rect -26 322 1074 521
rect -26 320 573 322
rect 47642 320 50758 519
<< obsm4 >>
rect -26 -328 50758 -320
<< metal5 >>
rect -26 900 692 1220
rect 47384 900 50758 1220
rect -26 260 692 580
rect 47704 579 50758 580
rect 47384 260 50758 579
<< obsm5 >>
rect -26 -328 50758 -320
use comparator  comparator_0
timestamp 1662929294
transform 1 0 23898 0 1 26079
box -1669 -1057 1961 897
use filter  filter_0
timestamp 1662974539
transform 1 0 1272 0 1 -2522
box -1298 2522 22766 33508
use filter  filter_1
timestamp 1662974539
transform -1 0 46804 0 1 -2522
box -1298 2522 22766 33508
use filter_clkgen  filter_clkgen_0
timestamp 1663630899
transform 1 0 20194 0 1 33977
box -1661 -2136 3360 1229
use level_shifter_low  level_shifter_low_0
timestamp 1663814281
transform 1 0 24311 0 1 33500
box -71 -46 2139 722
use level_shifter_low  level_shifter_low_1
timestamp 1663814281
transform 1 0 24311 0 -1 33504
box -71 -46 2139 722
use level_up_shifter_d_a  level_up_shifter_d_a_0
timestamp 1662953364
transform 1 0 8352 0 1 32786
box 402 498 2794 1683
use level_up_shifter_d_a  level_up_shifter_d_a_1
timestamp 1662953364
transform -1 0 39952 0 1 32786
box 402 498 2794 1683
<< labels >>
flabel metal2 37782 30236 37816 32872 1 FreeSans 1600 0 0 0 ctrl
flabel metal2 38301 30356 38335 32884 1 FreeSans 1600 0 0 0 ctrl_
flabel metal2 9969 33461 10003 33848 1 FreeSans 1600 0 0 0 fb
flabel metal2 10488 33460 10522 33848 1 FreeSans 1600 0 0 0 fb_inv
flabel metal2 5052 35140 5108 37140 1 FreeSans 1600 0 0 0 fb1
port 28 n default input
flabel metal2 13516 33032 13572 37140 1 FreeSans 1600 0 0 0 cclk
port 27 n default input
flabel metal2 21980 35470 22036 37140 1 FreeSans 1600 0 0 0 div2
port 29 n default input
flabel metal2 30444 35481 30500 37140 1 FreeSans 1600 0 0 0 high_buf
port 30 n default output
flabel metal2 38908 35457 38964 37140 1 FreeSans 1600 0 0 0 phi1b_dig
port 31 n default output
flabel metal2 47372 34983 47428 37140 1 FreeSans 1600 0 0 0 lo
port 32 n default input
<< end >>
