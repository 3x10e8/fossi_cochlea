magic
tech sky130A
magscale 1 2
timestamp 1647895372
<< nwell >>
rect -512 -6 1153 164
<< pwell >>
rect 2901 -332 2928 -210
rect 4626 -329 4659 -153
rect 6356 -332 6389 -156
rect 8075 -335 8108 -159
rect 8860 -276 8951 -200
rect 8860 -291 8871 -276
rect 8919 -303 8951 -276
rect 8846 -340 8894 -311
rect 8895 -358 8959 -305
rect 8891 -388 8959 -358
<< pmos >>
rect -418 34 -388 118
rect -330 34 -300 118
rect 0 34 30 118
rect 88 34 118 118
rect 176 34 206 118
rect 264 34 294 118
rect 528 30 558 114
rect 618 30 648 114
rect 902 30 932 114
rect 992 30 1022 114
<< nmoslvt >>
rect -430 -266 -400 -182
rect -324 -266 -294 -182
rect -104 -266 -74 -182
rect 0 -266 30 -182
rect 88 -266 118 -182
rect 176 -266 206 -182
rect 264 -266 294 -182
rect 528 -266 558 -182
rect 618 -266 648 -182
rect 902 -266 932 -182
rect 992 -266 1022 -182
<< ndiff >>
rect -504 -204 -430 -182
rect -504 -238 -496 -204
rect -462 -238 -430 -204
rect -504 -266 -430 -238
rect -400 -204 -324 -182
rect -400 -238 -378 -204
rect -344 -238 -324 -204
rect -400 -266 -324 -238
rect -294 -204 -220 -182
rect -294 -238 -262 -204
rect -228 -238 -220 -204
rect -294 -266 -220 -238
rect -158 -204 -104 -182
rect -158 -238 -150 -204
rect -116 -238 -104 -204
rect -158 -266 -104 -238
rect -74 -216 0 -182
rect -74 -250 -60 -216
rect -26 -250 0 -216
rect -74 -266 0 -250
rect 30 -204 88 -182
rect 30 -238 42 -204
rect 76 -238 88 -204
rect 30 -266 88 -238
rect 118 -204 176 -182
rect 118 -238 130 -204
rect 164 -238 176 -204
rect 118 -266 176 -238
rect 206 -204 264 -182
rect 206 -238 218 -204
rect 252 -238 264 -204
rect 206 -266 264 -238
rect 294 -204 354 -182
rect 294 -238 306 -204
rect 340 -238 354 -204
rect 294 -266 354 -238
rect 470 -204 528 -182
rect 470 -238 482 -204
rect 516 -238 528 -204
rect 470 -266 528 -238
rect 558 -204 618 -182
rect 558 -238 570 -204
rect 604 -238 618 -204
rect 558 -266 618 -238
rect 648 -204 708 -182
rect 648 -238 660 -204
rect 694 -238 708 -204
rect 842 -204 902 -182
rect 648 -266 708 -238
rect 842 -238 856 -204
rect 890 -238 902 -204
rect 842 -266 902 -238
rect 932 -204 992 -182
rect 932 -238 944 -204
rect 978 -238 992 -204
rect 932 -266 992 -238
rect 1022 -204 1080 -182
rect 1022 -238 1034 -204
rect 1068 -238 1080 -204
rect 1022 -266 1080 -238
<< pdiff >>
rect -476 96 -418 118
rect -476 62 -464 96
rect -430 62 -418 96
rect -476 34 -418 62
rect -388 96 -330 118
rect -388 62 -376 96
rect -342 62 -330 96
rect -388 34 -330 62
rect -300 96 -246 118
rect -300 62 -288 96
rect -254 62 -246 96
rect -300 34 -246 62
rect -54 96 0 118
rect -54 62 -46 96
rect -12 62 0 96
rect -54 34 0 62
rect 30 96 88 118
rect 30 62 42 96
rect 76 62 88 96
rect 30 34 88 62
rect 118 96 176 118
rect 118 62 130 96
rect 164 62 176 96
rect 118 34 176 62
rect 206 96 264 118
rect 206 62 218 96
rect 252 62 264 96
rect 206 34 264 62
rect 294 96 354 118
rect 294 62 306 96
rect 340 62 354 96
rect 294 34 354 62
rect 470 86 528 114
rect 470 52 482 86
rect 516 52 528 86
rect 470 30 528 52
rect 558 86 618 114
rect 558 52 572 86
rect 606 52 618 86
rect 558 30 618 52
rect 648 86 708 114
rect 648 52 660 86
rect 694 52 708 86
rect 842 86 902 114
rect 648 30 708 52
rect 842 52 856 86
rect 890 52 902 86
rect 842 30 902 52
rect 932 86 992 114
rect 932 52 946 86
rect 980 52 992 86
rect 932 30 992 52
rect 1022 86 1080 114
rect 1022 52 1034 86
rect 1068 52 1080 86
rect 1022 30 1080 52
<< ndiffc >>
rect -496 -238 -462 -204
rect -378 -238 -344 -204
rect -262 -238 -228 -204
rect -150 -238 -116 -204
rect -60 -250 -26 -216
rect 42 -238 76 -204
rect 130 -238 164 -204
rect 218 -238 252 -204
rect 306 -238 340 -204
rect 482 -238 516 -204
rect 570 -238 604 -204
rect 660 -238 694 -204
rect 856 -238 890 -204
rect 944 -238 978 -204
rect 1034 -238 1068 -204
<< pdiffc >>
rect -464 62 -430 96
rect -376 62 -342 96
rect -288 62 -254 96
rect -46 62 -12 96
rect 42 62 76 96
rect 130 62 164 96
rect 218 62 252 96
rect 306 62 340 96
rect 482 52 516 86
rect 572 52 606 86
rect 660 52 694 86
rect 856 52 890 86
rect 946 52 980 86
rect 1034 52 1068 86
<< psubdiff >>
rect 354 -206 416 -182
rect 354 -240 382 -206
rect 354 -266 416 -240
rect 708 -228 842 -182
rect 708 -262 770 -228
rect 804 -262 842 -228
rect 708 -266 842 -262
rect 8895 -312 8959 -305
rect 8847 -330 8959 -312
rect 8847 -364 8904 -330
rect 8946 -364 8959 -330
rect 8847 -372 8959 -364
rect 8891 -388 8959 -372
<< nsubdiff >>
rect 8826 265 8961 270
rect 8826 228 8871 265
rect 8909 228 8961 265
rect 8826 187 8961 228
rect 354 92 416 118
rect 354 58 382 92
rect 354 34 416 58
rect 708 110 842 114
rect 708 76 782 110
rect 816 76 842 110
rect 708 30 842 76
<< psubdiffcont >>
rect 382 -240 416 -206
rect 770 -262 804 -228
rect 8904 -364 8946 -330
<< nsubdiffcont >>
rect 8871 228 8909 265
rect 382 58 416 92
rect 782 76 816 110
<< poly >>
rect 150 230 216 246
rect 150 196 166 230
rect 200 226 216 230
rect 200 196 294 226
rect 150 186 216 196
rect -418 118 -388 144
rect -330 118 -300 144
rect 0 118 30 144
rect 88 118 118 144
rect 176 118 206 144
rect 264 118 294 196
rect -154 84 -70 100
rect -154 50 -144 84
rect -110 50 -70 84
rect -154 34 -70 50
rect 528 114 558 140
rect 618 114 648 140
rect 902 114 932 140
rect 992 114 1022 140
rect -418 14 -388 34
rect -330 14 -300 34
rect -418 -16 -204 14
rect -100 12 -70 34
rect 0 12 30 34
rect -246 -26 -172 -16
rect -100 -18 30 12
rect -246 -30 -170 -26
rect -236 -46 -170 -30
rect -204 -60 -170 -46
rect -204 -70 -100 -60
rect -446 -90 -382 -72
rect -446 -124 -432 -90
rect -398 -124 -382 -90
rect -446 -140 -382 -124
rect -340 -90 -278 -72
rect -340 -124 -326 -90
rect -292 -124 -278 -90
rect -340 -140 -278 -124
rect -204 -104 -152 -70
rect -118 -104 -100 -70
rect 88 -78 118 34
rect 176 2 206 34
rect 264 8 294 34
rect 168 -14 222 2
rect 168 -48 178 -14
rect 212 -48 222 -14
rect 168 -64 222 -48
rect 412 -36 466 -20
rect -204 -114 -100 -104
rect 72 -84 118 -78
rect 72 -100 126 -84
rect -430 -182 -400 -140
rect -324 -182 -294 -140
rect -430 -292 -400 -266
rect -324 -292 -294 -266
rect -204 -282 -174 -114
rect 72 -134 82 -100
rect 116 -134 126 -100
rect 72 -150 126 -134
rect -104 -182 -74 -156
rect 0 -182 30 -156
rect 88 -182 118 -150
rect 176 -182 206 -64
rect 412 -70 422 -36
rect 456 -38 466 -36
rect 528 -38 558 30
rect 456 -68 558 -38
rect 618 -58 648 30
rect 786 -36 840 -20
rect 456 -70 466 -68
rect 304 -94 358 -78
rect 412 -86 466 -70
rect 304 -114 314 -94
rect 264 -128 314 -114
rect 348 -128 358 -94
rect 264 -144 358 -128
rect 264 -182 294 -144
rect 528 -182 558 -68
rect 606 -74 660 -58
rect 606 -108 616 -74
rect 650 -108 660 -74
rect 786 -70 796 -36
rect 830 -38 840 -36
rect 902 -38 932 30
rect 830 -68 932 -38
rect 992 -58 1022 30
rect 830 -70 840 -68
rect 786 -86 840 -70
rect 606 -124 660 -108
rect 618 -182 648 -124
rect 902 -182 932 -68
rect 980 -74 1034 -58
rect 980 -108 990 -74
rect 1024 -108 1034 -74
rect 980 -124 1034 -108
rect 992 -182 1022 -124
rect -104 -282 -74 -266
rect -204 -312 -74 -282
rect 0 -334 30 -266
rect 88 -292 118 -266
rect 176 -292 206 -266
rect 264 -334 294 -266
rect 528 -292 558 -266
rect 618 -292 648 -266
rect 902 -292 932 -266
rect 992 -292 1022 -266
rect 0 -364 294 -334
<< polycont >>
rect 166 196 200 230
rect -144 50 -110 84
rect -432 -124 -398 -90
rect -326 -124 -292 -90
rect -152 -104 -118 -70
rect 178 -48 212 -14
rect 82 -134 116 -100
rect 422 -70 456 -36
rect 314 -128 348 -94
rect 616 -108 650 -74
rect 796 -70 830 -36
rect 990 -108 1024 -74
<< locali >>
rect -572 268 -510 302
rect -476 268 -414 302
rect -380 268 -318 302
rect -284 268 -222 302
rect -188 268 -126 302
rect -92 268 -30 302
rect 4 268 66 302
rect 100 268 162 302
rect 196 268 258 302
rect 292 268 354 302
rect 388 268 450 302
rect 484 268 546 302
rect 580 268 642 302
rect 676 268 738 302
rect 772 268 834 302
rect 868 268 930 302
rect 964 268 1026 302
rect 1060 268 1122 302
rect 1156 268 1218 302
rect -376 112 -342 268
rect -280 230 216 234
rect -280 200 166 230
rect -280 112 -246 200
rect 150 196 166 200
rect 200 196 216 230
rect 150 180 216 196
rect -504 96 -422 112
rect -504 62 -464 96
rect -430 62 -422 96
rect -504 46 -422 62
rect -384 96 -334 112
rect -384 62 -376 96
rect -342 62 -334 96
rect -384 46 -334 62
rect -296 110 -246 112
rect -296 96 -218 110
rect -296 62 -288 96
rect -254 62 -218 96
rect -296 46 -218 62
rect -504 -188 -470 46
rect -432 -90 -398 -72
rect -432 -140 -398 -124
rect -326 -90 -292 -72
rect -326 -140 -292 -124
rect -252 -188 -218 46
rect -150 84 -104 100
rect -150 50 -144 84
rect -110 50 -104 84
rect -150 34 -104 50
rect -54 96 -4 112
rect -54 62 -46 96
rect -12 62 -4 96
rect -54 46 -4 62
rect 34 96 84 112
rect 34 62 42 96
rect 76 62 84 96
rect 34 46 84 62
rect 122 96 176 112
rect 122 62 130 96
rect 164 62 176 96
rect 122 46 176 62
rect 210 96 260 112
rect 210 62 218 96
rect 252 62 260 96
rect 210 46 260 62
rect 298 96 348 112
rect 298 62 306 96
rect 340 62 348 96
rect 298 46 348 62
rect 382 92 416 268
rect 570 102 604 268
rect 782 110 816 268
rect -54 -14 -20 46
rect 178 -14 212 2
rect 306 -4 340 46
rect 382 42 416 58
rect 482 86 524 102
rect 516 52 524 86
rect 482 36 524 52
rect 564 86 614 102
rect 564 52 572 86
rect 606 52 614 86
rect 564 36 614 52
rect 652 86 736 102
rect 652 52 659 86
rect 694 52 736 86
rect 944 102 978 268
rect 782 60 816 76
rect 856 86 898 102
rect 652 36 736 52
rect 890 52 898 86
rect 856 36 898 52
rect 938 86 988 102
rect 938 52 946 86
rect 980 52 988 86
rect 938 36 988 52
rect 1026 86 1110 102
rect 1026 52 1034 86
rect 1068 52 1110 86
rect 1026 36 1110 52
rect -54 -48 178 -14
rect -168 -104 -152 -70
rect -118 -104 -102 -70
rect 14 -188 48 -48
rect 178 -64 212 -48
rect 246 -38 340 -4
rect 422 -36 456 -20
rect 82 -100 116 -84
rect 246 -100 280 -38
rect 116 -134 280 -100
rect 82 -150 116 -134
rect 220 -148 280 -134
rect 314 -94 348 -78
rect 422 -86 456 -70
rect 490 -74 524 36
rect 616 -74 650 -58
rect 314 -144 348 -128
rect 490 -108 616 -74
rect 220 -188 254 -148
rect 490 -188 524 -108
rect 616 -124 650 -108
rect 702 -188 736 36
rect 796 -36 830 -20
rect 796 -86 830 -70
rect 864 -74 898 36
rect 990 -74 1024 -58
rect 864 -108 990 -74
rect 864 -188 898 -108
rect 990 -124 1024 -108
rect 1076 -188 1110 36
rect 8354 -132 8392 -95
rect -504 -204 -454 -188
rect -504 -238 -496 -204
rect -462 -238 -454 -204
rect -504 -254 -454 -238
rect -386 -204 -336 -188
rect -386 -238 -378 -204
rect -344 -238 -336 -204
rect -386 -254 -336 -238
rect -270 -204 -218 -188
rect -270 -238 -262 -204
rect -228 -222 -218 -204
rect -156 -204 -108 -188
rect -228 -238 -220 -222
rect -270 -254 -220 -238
rect -156 -238 -150 -204
rect -116 -238 -108 -204
rect -156 -254 -108 -238
rect -66 -216 -20 -200
rect -66 -250 -60 -216
rect -26 -250 -20 -216
rect 14 -204 84 -188
rect 14 -222 42 -204
rect -380 -290 -346 -254
rect -156 -290 -122 -254
rect -66 -266 -20 -250
rect 34 -238 42 -222
rect 76 -238 84 -204
rect 34 -254 84 -238
rect 122 -204 172 -188
rect 122 -238 130 -204
rect 164 -238 172 -204
rect 122 -254 172 -238
rect 210 -204 260 -188
rect 210 -238 218 -204
rect 252 -238 260 -204
rect 210 -254 260 -238
rect 298 -204 348 -188
rect 298 -238 306 -204
rect 340 -238 348 -204
rect 298 -254 348 -238
rect 382 -206 416 -188
rect -380 -324 -122 -290
rect -54 -364 -20 -266
rect 132 -364 166 -254
rect 308 -364 342 -254
rect 382 -364 416 -240
rect 482 -204 524 -188
rect 516 -238 524 -204
rect 482 -254 524 -238
rect 562 -204 612 -188
rect 562 -238 570 -204
rect 604 -238 612 -204
rect 562 -254 612 -238
rect 652 -204 736 -188
rect 652 -238 660 -204
rect 694 -238 736 -204
rect 856 -204 898 -188
rect 652 -254 736 -238
rect 770 -228 804 -212
rect 572 -364 606 -254
rect 890 -238 898 -204
rect 856 -254 898 -238
rect 936 -204 986 -188
rect 936 -238 944 -204
rect 978 -238 986 -204
rect 936 -254 986 -238
rect 1026 -204 1110 -188
rect 1026 -238 1034 -204
rect 1068 -238 1110 -204
rect 1026 -254 1110 -238
rect 770 -364 804 -262
rect 946 -364 980 -254
rect 8904 -330 8946 -311
rect -572 -398 -510 -364
rect -476 -398 -414 -364
rect -380 -398 -318 -364
rect -284 -398 -222 -364
rect -188 -398 -126 -364
rect -92 -398 -30 -364
rect 4 -398 66 -364
rect 100 -398 162 -364
rect 196 -398 258 -364
rect 292 -398 354 -364
rect 388 -398 450 -364
rect 484 -398 546 -364
rect 580 -398 642 -364
rect 676 -398 738 -364
rect 772 -398 834 -364
rect 868 -398 930 -364
rect 964 -398 1026 -364
rect 1060 -398 1122 -364
rect 1156 -398 1218 -364
rect 8904 -372 8946 -364
<< viali >>
rect -510 268 -476 302
rect -414 268 -380 302
rect -318 268 -284 302
rect -222 268 -188 302
rect -126 268 -92 302
rect -30 268 4 302
rect 66 268 100 302
rect 162 268 196 302
rect 258 268 292 302
rect 354 268 388 302
rect 450 268 484 302
rect 546 268 580 302
rect 642 268 676 302
rect 738 268 772 302
rect 834 268 868 302
rect 930 268 964 302
rect 1026 268 1060 302
rect 1122 268 1156 302
rect -464 62 -430 96
rect -432 -124 -398 -90
rect -326 -124 -292 -90
rect -144 50 -110 84
rect 130 62 164 96
rect 659 52 660 86
rect 660 52 694 86
rect 4482 86 4516 120
rect 9182 91 9216 125
rect 178 -48 212 -14
rect -152 -104 -118 -70
rect 422 -70 456 -36
rect 82 -134 116 -100
rect 314 -128 348 -94
rect 796 -70 830 -36
rect 2754 5 2788 39
rect 6212 -17 6246 17
rect 8616 -6 8650 28
rect 3319 -71 3353 -37
rect 5047 -71 5081 -37
rect 6775 -71 6809 -37
rect 1234 -129 1268 -95
rect 1591 -117 1627 -79
rect 2962 -129 2996 -95
rect 4690 -129 4724 -95
rect 6418 -129 6452 -95
rect 7936 -132 7974 -95
rect 8135 -124 8175 -90
rect 8310 -111 8344 -77
rect 8826 -81 8862 -45
rect 9001 -75 9039 -41
rect 9293 -141 9329 -103
rect 8523 -186 8557 -152
rect 9470 -226 9506 -188
rect -510 -398 -476 -364
rect -414 -398 -380 -364
rect -318 -398 -284 -364
rect -222 -398 -188 -364
rect -126 -398 -92 -364
rect -30 -398 4 -364
rect 66 -398 100 -364
rect 162 -398 196 -364
rect 258 -398 292 -364
rect 354 -398 388 -364
rect 450 -398 484 -364
rect 546 -398 580 -364
rect 642 -398 676 -364
rect 738 -398 772 -364
rect 834 -398 868 -364
rect 930 -398 964 -364
rect 1026 -398 1060 -364
rect 1122 -398 1156 -364
<< metal1 >>
rect -572 302 1218 334
rect -572 268 -510 302
rect -476 268 -414 302
rect -380 268 -318 302
rect -284 268 -222 302
rect -188 268 -126 302
rect -92 268 -30 302
rect 4 268 66 302
rect 100 268 162 302
rect 196 268 258 302
rect 292 268 354 302
rect 388 268 450 302
rect 484 268 546 302
rect 580 268 642 302
rect 676 268 738 302
rect 772 268 834 302
rect 868 268 930 302
rect 964 268 1026 302
rect 1060 268 1122 302
rect 1156 268 1218 302
rect -572 236 1218 268
rect -476 98 -422 104
rect 130 102 164 236
rect 4470 120 4528 132
rect -476 96 -104 98
rect -476 62 -464 96
rect -430 84 -104 96
rect -430 62 -144 84
rect -476 60 -144 62
rect -476 54 -422 60
rect -150 50 -144 60
rect -110 50 -104 84
rect 124 96 170 102
rect 124 62 130 96
rect 164 62 170 96
rect 124 50 170 62
rect 648 86 707 100
rect 4470 86 4482 120
rect 4516 117 4528 120
rect 9169 125 9232 137
rect 5035 117 8322 119
rect 4516 86 8322 117
rect 648 52 659 86
rect 694 52 1629 86
rect 4470 85 8322 86
rect 4470 74 4528 85
rect -150 36 -104 50
rect 648 39 707 52
rect 168 -14 222 2
rect 168 -48 178 -14
rect 212 -36 466 -14
rect 212 -48 422 -36
rect -450 -72 -398 -69
rect -325 -71 -249 -65
rect -450 -78 -382 -72
rect -398 -130 -382 -78
rect -450 -140 -382 -130
rect -340 -79 -249 -71
rect -340 -131 -326 -79
rect -274 -131 -249 -79
rect -175 -115 -168 -58
rect -107 -115 -96 -58
rect 168 -64 222 -48
rect 412 -70 422 -48
rect 456 -70 466 -36
rect 72 -100 126 -82
rect -340 -140 -249 -131
rect -450 -143 -398 -140
rect -325 -147 -249 -140
rect 72 -134 82 -100
rect 116 -134 126 -100
rect 72 -150 126 -134
rect 305 -83 360 -76
rect 305 -136 308 -83
rect 412 -86 466 -70
rect 790 -36 840 -14
rect 790 -70 796 -36
rect 830 -70 840 -36
rect 1591 -70 1629 52
rect 2742 39 2801 46
rect 2742 5 2754 39
rect 2788 5 3369 39
rect 2742 -3 2801 5
rect 3304 -37 3369 5
rect 5046 -27 5089 85
rect 6199 17 6260 29
rect 6199 -17 6212 17
rect 6246 -17 6815 17
rect 790 -86 840 -70
rect 1222 -83 1280 -77
rect 305 -147 360 -136
rect 82 -204 116 -150
rect 796 -204 830 -86
rect 1580 -79 1637 -70
rect 3304 -71 3319 -37
rect 3353 -71 3369 -37
rect 1580 -117 1591 -79
rect 1627 -117 1637 -79
rect 1580 -125 1637 -117
rect 2940 -85 3021 -71
rect 3304 -77 3369 -71
rect 5035 -37 5095 -27
rect 6199 -29 6260 -17
rect 5035 -71 5047 -37
rect 5081 -71 5095 -37
rect 1591 -139 1629 -125
rect 2940 -137 2955 -85
rect 3007 -137 3021 -85
rect 1222 -147 1280 -141
rect 2940 -152 3021 -137
rect 4671 -85 4748 -72
rect 5035 -78 5095 -71
rect 6763 -37 6815 -17
rect 6763 -71 6775 -37
rect 6809 -71 6815 -37
rect 8285 -60 8322 85
rect 9169 91 9182 125
rect 9216 91 9624 125
rect 9169 79 9232 91
rect 8603 28 9054 37
rect 8603 -6 8616 28
rect 8650 -1 9054 28
rect 8650 -6 8666 -1
rect 8603 -12 8666 -6
rect 8788 -45 8933 -32
rect 4671 -137 4683 -85
rect 4735 -137 4748 -85
rect 4671 -151 4748 -137
rect 6394 -85 6475 -74
rect 6394 -138 6409 -85
rect 6461 -138 6475 -85
rect 6763 -97 6815 -71
rect 8255 -62 8443 -60
rect 8788 -62 8826 -45
rect 8255 -77 8826 -62
rect 7930 -90 8189 -81
rect 7930 -95 8135 -90
rect 6394 -153 6475 -138
rect 7930 -132 7936 -95
rect 7974 -124 8135 -95
rect 8175 -124 8189 -90
rect 7974 -132 8189 -124
rect 8255 -111 8310 -77
rect 8344 -81 8826 -77
rect 8862 -81 8933 -45
rect 8344 -111 8933 -81
rect 8979 -41 9054 -1
rect 8979 -75 9001 -41
rect 9039 -75 9054 -41
rect 8979 -83 9054 -75
rect 9281 -103 9341 -86
rect 8255 -127 8443 -111
rect 7930 -146 8189 -132
rect 9281 -141 9293 -103
rect 9329 -141 9341 -103
rect 8509 -150 8571 -141
rect 9281 -150 9341 -141
rect 8509 -152 9341 -150
rect 8509 -186 8523 -152
rect 8557 -186 9341 -152
rect 8509 -200 8571 -186
rect 9458 -188 9518 -176
rect 82 -238 830 -204
rect 9458 -226 9470 -188
rect 9506 -190 9518 -188
rect 9506 -224 9642 -190
rect 9506 -226 9518 -224
rect 9458 -239 9518 -226
rect -572 -364 1218 -332
rect -572 -398 -510 -364
rect -476 -398 -414 -364
rect -380 -398 -318 -364
rect -284 -398 -222 -364
rect -188 -398 -126 -364
rect -92 -398 -30 -364
rect 4 -398 66 -364
rect 100 -398 162 -364
rect 196 -398 258 -364
rect 292 -398 354 -364
rect 388 -398 450 -364
rect 484 -398 546 -364
rect 580 -398 642 -364
rect 676 -398 738 -364
rect 772 -398 834 -364
rect 868 -398 930 -364
rect 964 -398 1026 -364
rect 1060 -398 1122 -364
rect 1156 -398 1218 -364
rect -572 -430 1218 -398
<< via1 >>
rect -450 -90 -398 -78
rect -450 -124 -432 -90
rect -432 -124 -398 -90
rect -450 -130 -398 -124
rect -326 -90 -274 -79
rect -326 -124 -292 -90
rect -292 -124 -274 -90
rect -326 -131 -274 -124
rect -168 -70 -107 -58
rect -168 -104 -152 -70
rect -152 -104 -118 -70
rect -118 -104 -107 -70
rect -168 -115 -107 -104
rect 308 -94 360 -83
rect 308 -128 314 -94
rect 314 -128 348 -94
rect 348 -128 360 -94
rect 308 -136 360 -128
rect 1222 -95 1280 -83
rect 1222 -129 1234 -95
rect 1234 -129 1268 -95
rect 1268 -129 1280 -95
rect 1222 -141 1280 -129
rect 2955 -95 3007 -85
rect 2955 -129 2962 -95
rect 2962 -129 2996 -95
rect 2996 -129 3007 -95
rect 2955 -137 3007 -129
rect 4683 -95 4735 -85
rect 4683 -129 4690 -95
rect 4690 -129 4724 -95
rect 4724 -129 4735 -95
rect 4683 -137 4735 -129
rect 6409 -95 6461 -85
rect 6409 -129 6418 -95
rect 6418 -129 6452 -95
rect 6452 -129 6461 -95
rect 6409 -138 6461 -129
<< metal2 >>
rect -574 30 -544 401
rect -364 219 -334 374
rect -364 189 338 219
rect -574 1 -99 30
rect -146 -58 -99 1
rect -464 -76 -398 -67
rect -325 -73 -249 -65
rect -407 -78 -398 -76
rect -407 -138 -398 -130
rect -326 -74 -249 -73
rect -326 -79 -315 -74
rect -326 -137 -315 -131
rect -464 -147 -398 -138
rect -325 -138 -315 -137
rect -259 -138 -249 -74
rect -175 -115 -168 -58
rect -107 -115 -96 -58
rect 305 -72 338 189
rect 304 -81 363 -72
rect -325 -147 -249 -138
rect 304 -139 306 -81
rect 362 -139 363 -81
rect 304 -148 363 -139
rect 1216 -77 1289 -68
rect 1216 -147 1222 -77
rect 1280 -147 1289 -77
rect 1216 -156 1289 -147
rect 2940 -80 3021 -71
rect 2940 -143 2949 -80
rect 3012 -143 3021 -80
rect 2940 -152 3021 -143
rect 4671 -81 4748 -72
rect 4671 -142 4680 -81
rect 4739 -142 4748 -81
rect 4671 -151 4748 -142
rect 6394 -84 6475 -74
rect 6394 -144 6404 -84
rect 6465 -144 6475 -84
rect 6394 -153 6475 -144
<< via2 >>
rect -464 -78 -407 -76
rect -464 -130 -450 -78
rect -450 -130 -407 -78
rect -464 -138 -407 -130
rect -315 -79 -259 -74
rect -315 -131 -274 -79
rect -274 -131 -259 -79
rect -315 -138 -259 -131
rect 306 -83 362 -81
rect 306 -136 308 -83
rect 308 -136 360 -83
rect 360 -136 362 -83
rect 306 -139 362 -136
rect 1222 -83 1280 -77
rect 1222 -141 1280 -83
rect 1222 -147 1280 -141
rect 2949 -85 3012 -80
rect 2949 -137 2955 -85
rect 2955 -137 3007 -85
rect 3007 -137 3012 -85
rect 2949 -143 3012 -137
rect 4680 -85 4739 -81
rect 4680 -137 4683 -85
rect 4683 -137 4735 -85
rect 4735 -137 4739 -85
rect 4680 -142 4739 -137
rect 6404 -85 6465 -84
rect 6404 -138 6409 -85
rect 6409 -138 6461 -85
rect 6461 -138 6465 -85
rect 6404 -144 6465 -138
<< metal3 >>
rect -555 -73 -398 -69
rect -555 -140 -472 -73
rect -407 -140 -398 -73
rect -555 -144 -398 -140
rect -326 -72 -169 -69
rect -326 -139 -315 -72
rect -251 -139 -169 -72
rect -326 -144 -169 -139
rect 300 -81 367 -72
rect 1216 -77 1289 -68
rect 1216 -79 1222 -77
rect 1173 -81 1222 -79
rect 300 -139 306 -81
rect 362 -139 1222 -81
rect 300 -146 1222 -139
rect 300 -148 367 -146
rect 1216 -147 1222 -146
rect 1280 -79 1289 -77
rect 2940 -79 3021 -71
rect 4671 -79 4748 -72
rect 6394 -79 6475 -74
rect 1280 -80 6475 -79
rect 1280 -143 2949 -80
rect 3012 -81 6475 -80
rect 3012 -142 4680 -81
rect 4739 -84 6475 -81
rect 4739 -142 6404 -84
rect 3012 -143 6404 -142
rect 1280 -144 6404 -143
rect 6465 -144 6475 -84
rect 1280 -146 6475 -144
rect 1280 -147 1289 -146
rect 1216 -156 1289 -147
rect 2940 -152 3021 -146
rect 4671 -151 4748 -146
rect 6394 -153 6475 -146
<< via3 >>
rect -472 -76 -407 -73
rect -472 -138 -464 -76
rect -464 -138 -407 -76
rect -472 -140 -407 -138
rect -315 -74 -251 -72
rect -315 -138 -259 -74
rect -259 -138 -251 -74
rect -315 -139 -251 -138
<< metal4 >>
rect -274 -69 -196 -42
rect -476 -73 -404 -71
rect -476 -74 -472 -73
rect -555 -134 -472 -74
rect -476 -140 -472 -134
rect -407 -140 -404 -73
rect -476 -142 -404 -140
rect -318 -72 -196 -69
rect -318 -139 -315 -72
rect -251 -139 -196 -72
rect -318 -141 -196 -139
use sky130_fd_sc_lp__buf_1  sky130_fd_sc_lp__buf_1_0 /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1647888116
transform -1 0 9539 0 1 -381
box -38 -49 326 715
use sky130_fd_sc_lp__and2_1  sky130_fd_sc_lp__and2_1_0 /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1626515395
transform 1 0 8771 0 1 -381
box -38 -49 518 715
use sky130_fd_sc_lp__xor2_1  sky130_fd_sc_lp__xor2_1_0 /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1640850677
transform 1 0 8099 0 1 -381
box -38 -49 710 715
use sky130_fd_sc_lp__dfxtp_2  sky130_fd_sc_lp__dfxtp_2_0 /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_lp/mag
timestamp 1647887894
transform 1 0 1187 0 1 -381
box -38 -49 1766 715
use sky130_fd_sc_lp__dfxtp_2  sky130_fd_sc_lp__dfxtp_2_1
timestamp 1647887894
transform 1 0 2915 0 1 -381
box -38 -49 1766 715
use sky130_fd_sc_lp__dfxtp_2  sky130_fd_sc_lp__dfxtp_2_2
timestamp 1647887894
transform 1 0 4643 0 1 -381
box -38 -49 1766 715
use sky130_fd_sc_lp__dfxtp_2  sky130_fd_sc_lp__dfxtp_2_3
timestamp 1647887894
transform 1 0 6371 0 1 -381
box -38 -49 1766 715
<< labels >>
flabel polycont 178 -48 212 -14 0 FreeSans 112 0 0 0 high
flabel polycont 82 -134 116 -100 0 FreeSans 112 0 0 0 low
flabel polycont 314 -128 348 -94 0 FreeSans 112 0 0 0 phi1b
flabel polycont -152 -104 -118 -70 0 FreeSans 112 0 0 0 phi1
rlabel locali -102 -88 -102 -88 3 phi1
rlabel locali 236 112 236 112 1 pfete
rlabel locali 60 112 60 112 1 pfetw
rlabel locali 236 -188 236 -188 1 low
rlabel locali 60 -188 60 -188 1 high
rlabel locali 330 -78 330 -78 1 phi1b
rlabel locali -208 -290 -208 -290 1 tail
rlabel locali -310 -74 -310 -74 1 inm
flabel polycont -326 -124 -292 -90 0 FreeSans 112 0 0 0 inm
flabel polycont -432 -124 -398 -90 0 FreeSans 112 0 0 0 inp
rlabel locali -414 -72 -414 -72 1 inp
rlabel locali -470 -40 -470 -40 3 FP
rlabel locali -252 -46 -252 -46 7 FN
rlabel locali 546 288 546 288 3 VDD
rlabel locali 546 -382 546 -382 3 GND
flabel pdiffc 660 52 694 86 0 FreeSans 112 0 0 0 high_buffered
flabel ndiffc 1034 -238 1068 -204 0 FreeSans 112 0 0 0 low_buffered
flabel space 1539 -71 1754 -34 0 FreeSans 160 0 0 0 compout
flabel space 3291 -53 3506 -16 0 FreeSans 160 0 0 0 latch
flabel space 4971 -29 5186 8 0 FreeSans 160 0 0 0 pol_1
flabel space 7863 107 8078 144 0 FreeSans 160 0 0 0 pol_2
rlabel metal1 9642 -207 9642 -207 3 events
rlabel metal1 9624 107 9624 107 3 polxevent
flabel space 9324 -316 9536 -124 0 FreeSans 800 0 0 0 Events
flabel space 9110 77 9547 155 0 FreeSans 480 0 0 0 polxevent
<< end >>
